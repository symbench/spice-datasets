.title KiCad schematic
N2 20190121
N1 OHWLOGO
J3 GND NC_01 /POWER_0 Conn_01x03
J4 GND NC_02 /POWER_1 Conn_01x03
J5 /POWER_0 GND /POWER_1 GND /SIGNAL_0 Net-_J5-Pad6_ /SIGNAL_1 Net-_J5-Pad8_ /SIGNAL_2 Net-_J5-Pad10_ Conn_02x05_Odd_Even
C1 /POWER_0 GND C
C2 /POWER_1 GND C
R4 /SIGNAL_0 /SIGNAL R
R7 GND /SIGNAL_0 R
R1 GND /SIGNAL R
R5 /SIGNAL_1 /SIGNAL R
R8 GND /SIGNAL_1 R
R2 GND /SIGNAL R
R6 /SIGNAL_2 /SIGNAL R
R9 GND /SIGNAL_2 R
R3 GND /SIGNAL R
J1 GND /SIGNAL Coax
SJ1 Net-_J5-Pad6_ GND SolderJumper_2way_1conn
SJ2 Net-_J5-Pad8_ GND SolderJumper_2way_1conn
SJ3 Net-_J5-Pad10_ GND SolderJumper_2way_1conn
.end
