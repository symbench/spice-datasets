.title KiCad schematic
U5 NC_01 NC_02 NC_03 Net-_U5-Pad5_ Net-_U5-Pad6_ NC_04 NC_05 NC_06 NC_07 /TIM2_CH1 /TIM2_CH2 /rot_but NC_08 NC_09 /ADC1_IN5 /ADC1_IN6 /ADC1_IN7 NC_10 NC_11 NC_12 NC_13 BOOT /DISP_SCL /I2S2_WS /I2S2_CK /I2S2ext /I2S2_SD /I2S2_MCK NC_14 /SDIO_D0 /SDIO_D1 NC_15 /USART1_TX /USART1_RX /stomp_start /stomp_stop Net-_J3-Pad4_ Net-_J3-Pad2_ /SDdetect /SDIO_D2 /SDIO_D3 /SDIO_CK /SDIO_CMD /DISP_SDA NC_16 NC_17 /I2C1_SCL /I2C1_SDA NC_18 NC_19 STM32F401RC
J3 3.3V Net-_J3-Pad2_ GND Net-_J3-Pad4_ programming header
U1 NC_20 NC_21 /I2S2_CK /I2S2_MCK /I2S2_SD /I2S2_WS /I2S2_CK /I2S2_MCK /I2S2ext /I2S2_WS GND GND /I2C1_SDA /I2C1_SCL WM8778-units
SW2 GND BOOT 3.3V RAM~FLASH
J4 /SDIO_D2 /SDIO_D3 /SDIO_CMD 3.3V /SDIO_CK GND /SDIO_D0 /SDIO_D1 GND /SDdetect GND Micro_SD_Card_Det
R6 3.3V /I2C1_SDA 4.7k
R5 3.3V /I2C1_SCL 4.7k
R4 3.3V /SDdetect 4.7k
SW5 /TIM2_CH2 /TIM2_CH1 GND /rot_but GND Rotary_Encoder_Switch
R7 /rot_but 3.3V 4.7k
C33 /rot_but GND 100nF
U6 GND 3.3V /DISP_SCL /DISP_SDA lcd
RV1 GND /ADC1_IN5 3.3V pot_in_l
RV2 GND /ADC1_IN6 3.3V pot_in_r
RV3 GND /ADC1_IN7 3.3V pot_out
SW3 /stomp_start GND start
SW4 /stomp_stop GND stop
J2 /USART1_RX /USART1_TX UART
C32 GND 3.3V 10uF
C31 GND 3.3V 4.7uF
Y1 Net-_U5-Pad5_ GND Net-_U5-Pad6_ CSTLS4M00G53-B0
.end
