.title KiCad schematic
U1 NC_01 NC_02 NC_03 +5V GND NC_04 Net-_C4-Pad1_ Net-_C3-Pad1_ NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 SpdMOSI SpdMISO SpdSCK +5V NC_11 Net-_C1-Pad1_ GND NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 SpdRESET SpdRXD SpdTXD NC_19 ATmega328PB-AU
Y1 Net-_C3-Pad1_ Net-_C4-Pad1_ Crystal
C3 Net-_C3-Pad1_ GND C
C4 Net-_C4-Pad1_ GND C
C5 +5V GND C
C1 Net-_C1-Pad1_ GND C
D1 Net-_C1-Pad1_ GND LM4040DBZ-3
R1 +5V Net-_C1-Pad1_ R
R2 +5V SpdRESET R
C2 SpdRESET GND C
J1 SpdMISO +5V SpdSCK SpdMOSI SpdRESET GND AVR-ISP-6
J2 SpdDTR SpdTXD SpdRXD +5V GND GND FTDI_Header
C6 SpdRESET SpdDTR C
.end
