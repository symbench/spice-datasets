.title KiCad schematic
J1 /Vcc /GND /12V /9V /5V /3.3V Conn_01x06
J2 Net-_J2-Pad1_ Net-_J2-Pad2_ Conn_01x02
T1 Net-_J2-Pad2_ Net-_J2-Pad1_ Net-_D1-Pad4_ Net-_D1-Pad3_ Transformer_1P_1S
D1 /Vcc /GND Net-_D1-Pad3_ Net-_D1-Pad4_ FB_RECT
C1 /Vcc /GND 470uF 50v
U1 Net-_C2-Pad1_ NC_01 NC_02 /12V Net-_R1-Pad2_ /GND /Vcc Net-_C2-Pad2_ LM2675M-12
R1 /Vcc Net-_R1-Pad2_ 10k
D2 Net-_C2-Pad2_ /GND D_Schottky
C3 /12V /GND CP1_Small
L1 Net-_C2-Pad2_ /12V 47uH
C2 Net-_C2-Pad1_ Net-_C2-Pad2_ 10nF
R2 /Vcc Net-_R2-Pad2_ 10k
D3 Net-_C4-Pad2_ /GND D_Schottky
C5 /9V /GND CP1_Small
L2 Net-_C4-Pad2_ /9V 47uH
C4 Net-_C4-Pad1_ Net-_C4-Pad2_ 10nF
R4 /9V Net-_R3-Pad2_ 9.1k
R3 /GND Net-_R3-Pad2_ 1.4k
U2 Net-_C4-Pad1_ NC_03 NC_04 Net-_R3-Pad2_ Net-_R2-Pad2_ /GND /Vcc Net-_C4-Pad2_ LM2675M-ADJ
R5 /Vcc Net-_R5-Pad2_ 10k
D4 Net-_C6-Pad2_ /GND D_Schottky
C7 /5V /GND CP1_Small
L3 Net-_C6-Pad2_ /5V 47uH
C6 Net-_C6-Pad1_ Net-_C6-Pad2_ 10nF
U3 Net-_C6-Pad1_ NC_05 NC_06 /5V Net-_R5-Pad2_ /GND /Vcc Net-_C6-Pad2_ LM2675M-5
R6 /Vcc Net-_R6-Pad2_ 10k
D5 Net-_C8-Pad2_ /GND D_Schottky
C9 /3.3V /GND CP1_Small
L4 Net-_C8-Pad2_ /3.3V 47uH
C8 Net-_C8-Pad1_ Net-_C8-Pad2_ 10nF
U4 Net-_C8-Pad1_ NC_07 NC_08 /3.3V Net-_R6-Pad2_ /GND /Vcc Net-_C8-Pad2_ LM2675M-3.3
.end
