.title KiCad schematic
U1 NC_01 NC_02 NC_03 NC_04 Net-_R1-Pad1_ NC_05 Net-_R2-Pad1_ NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 GND FPGA_Pluto
R1 Net-_R1-Pad1_ Measure_at_the_scope 47k
R2 Net-_R2-Pad1_ Measure_at_the_scope 1k
C1 Measure_at_the_scope GND 10n
.end
