.title KiCad schematic
P1 /5V /PWR_IO /3V3 CONN_01X03
R1 /DEVICE_RX /TEENCY_TX R
R2 /TEENCY_RX /DEVICE_TX R
U1 /TEENCY_RX /TEENCY_TX NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 /SPI_CS /SPI_MOSI /SPI_MISO /SPI_CLK /AIO_0 /AIO_1 /AIO_2 /AIO_3 /I2C_DAT /I2C_SCLK NC_09 NC_10 NC_11 NC_12 /3V3 NC_13 /5V /GND NC_14 NC_15 /GND NC_16 NC_17 Teensy-3.2
H1 /PWR_IO /SPI_MOSI /SPI_MISO /SPI_CLK /SPI_CS /DEVICE_RX /DEVICE_TX /GND /3V3 /I2C_SCLK /I2C_DAT /AIO_0 /AIO_1 /AIO_2 /AIO_3 /GND CE_Header
R3 /I2C_SCLK /3V3 4.7kΩ
R4 /I2C_DAT /3V3 4.7kΩ
.end
