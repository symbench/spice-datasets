.title KiCad schematic
U14 NC_01 NC_02 GND GND GND /TX_ISOLATED /RX_ISOLATED /GPS_VCC /GPS_VCC /GPS_VCC NC_03 NC_04 MAX-M8Q
U13 /RX_ISOLATED GND +3V3 NC_05 NC_06 /GPS_VCC /GPS_VCC /TX_ISOLATED TXB0102DCU
C52 +3V3 GND 0.1uF
R29 /GPS_VCC GND 100K
U15 +3V3 GND CC_GPIO8 Net-_C59-Pad1_ /GPS_VCC /GPS_VCC TPS22918
C59 Net-_C59-Pad1_ GND 0.001uF
R32 CC_GPIO8 GND 100K
C61 GND +3V3 1uF
C57 /GPS_VCC GND 22uF
.end
