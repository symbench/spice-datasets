.title KiCad schematic
D1 NC_01 NC_02 NC_03 NC_04 Diode_Bridge
.end
