.title KiCad schematic
U1 /!MCLR NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 +5V GND NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 GND +5V NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 PIC18F452-IP
Y1 NC_36 NC_37 Crystal
R1 +5V Net-_C1-Pad1_ 10K
C1 Net-_C1-Pad1_ GND C
R2 /!MCLR Net-_C1-Pad1_ 510
SW1 NC_38 Net-_C1-Pad1_ NC_39 GND SW_Push_Dual
.end
