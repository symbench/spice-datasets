.title KiCad schematic
J2 GND NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NEIGHBOR2
J1 GND VCC NC_40 /P0_0 NC_41 /P0_1 NC_42 NC_43 NC_44 NC_45 NC_46 NC_47 NC_48 NC_49 NC_50 NC_51 NC_52 NC_53 NC_54 NC_55 NC_56 NC_57 NC_58 NC_59 NC_60 NC_61 NC_62 NC_63 NC_64 NC_65 NC_66 NC_67 NC_68 NC_69 NC_70 NC_71 NC_72 NC_73 NC_74 NC_75 NEIGHBOR1
J7 GND NC_76 NC_77 NC_78 NC_79 NC_80 NC_81 NC_82 NC_83 GND NC_84 NC_85 NC_86 NC_87 NC_88 NC_89 NC_90 NC_91 GND NC_92 BONUS_ROW
MH3 GND MOUNTING_HOLE
MH4 GND MOUNTING_HOLE
MH1 GND MOUNTING_HOLE
MH2 GND MOUNTING_HOLE
U1 /+IN_A /-IN_A /+IN_B /-IN_B GND /OUT_B /OUT_A VCC TLV3502
C1 GND VCC C
R14 /-IN_A GND R
R16 /+IN_A GND R
R10 /-IN_B GND R
R12 /+IN_B GND R
R13 VCC /-IN_A R
R15 VCC /+IN_A R
R9 VCC /-IN_B R
R11 VCC /+IN_B R
R3 /+IN_A /RXBBQ- 0
R4 /-IN_A /RXBBQ+ 0
R5 /+IN_B /RXBBI- 0
R6 /-IN_B /RXBBI+ 0
R7 /+IN_A /-IN_A R
R8 /+IN_B /-IN_B R
P9 GND GND GND /RXBBQ- /RXBBI- /RXBBQ+ /RXBBI+ GND GND NC_93 NC_94 NC_95 NC_96 GND GND GND BASEBAND
R1 /P0_1 /OUT_A 0
R2 /P0_0 /OUT_B 0
.end
