.title KiCad schematic
U1 NC_01 HOLE
U2 NC_02 HOLE
U3 NC_03 HOLE
U4 NC_04 HOLE
U5 +5V +3V3 NC_05 NC_06 NC_07 NC_08 /A4 /A5 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 GND GND GND IOREF NC_24 NC_25 /A5 /A4 VIN ARDUINO-101-SHIELD
.end
