.title KiCad schematic
U1 /G2 /INT /OUT /BIAS VCC /IN+ /IN- GND /AUX_IN /G1 MAX4062
R3 /G1 /G2 11K
C6 Net-_C6-Pad1_ /IN+ 1uf
C5 GND /IN- 1uf
C4 Net-_C4-Pad1_ /AUX_IN 1uf
C7 VCC GND 100n
C1 GND /BIAS 100n
R2 /INT VCC 100K
J3 GND /OUT OUT
J4 GND Net-_C4-Pad1_ AUX
J5 GND Net-_C6-Pad1_ MIC
J1 GND +9V PWR
J2 Net-_J2-Pad1_ INT
R1 /INT Net-_J2-Pad1_ 100
U2 +9V +9V +9V NC_01 GND +9V Net-_C3-Pad1_ GND VCC VCC LT3042
R4 GND Net-_C3-Pad1_ 50K
C2 +9V GND 10uf
C8 VCC GND 10uf
C3 Net-_C3-Pad1_ GND 0.47uf
.end
