.title KiCad schematic
J14 eDP_VCC eDP_VCC GSENS_VCC TOUCH_VCC CAM_P_1 CAM_VCC NC_01 NC_02 NC_03 GND NC_04 NC_05 GND NC_06 NC_07 GND NC_08 NC_09 GND NC_10 NC_11 TOUCH_P_1 TOUCH_D1 TOUCH_D2 GND NC_12 NC_13 GND NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 eDP_VLED eDP_VLED eDP_VLED GND LENOVO_FPC
J1 NC_23 NC_24 NC_25 NC_26 GND GND CAM_U
J4 NC_27 NC_28 NC_29 GND GND MIC_S
J7 NC_30 NC_31 NC_32 GND MIC
J3 NC_33 NC_34 CAM_EN
J8 CAM_VCC GND CAM_VCC
J9 GSENS_VCC NC_35 NC_36 NC_37 GND GSENS_PI
J5 NC_38 NC_39 NC_40 NC_41 GND GSENS_S
J2 NC_42 TOUCH_D2 TOUCH_D1 NC_43 GND GND TOUCH_U
J13 TOUCH_VCC TOUCH_D1 TOUCH_D2 GND GND TOUCH_S
J6 TOUCH_P_1 GND TOUCH_P1
J11 TOUCH_VCC GND TOUCH_VCC
J12 TOUCH_VCC TOUCH_D1 TOUCH_D2 TOUCH_P_1 GND TOUCH
J10 CAM_VCC NC_44 NC_45 CAM_P_1 GND CAM
J15 NC_46 NC_47 NC_48 NC_49 NC_50 CAM_S
.end
