.title KiCad schematic
U1 GNDA Net-_R1-Pad2_ Net-_C17-Pad1_ GNDA Net-_C4-Pad1_ VDD VSS xStby xMute VDD /OutL VSS TDA7294V
C7 GND VSS 220n
C8 GND VSS 2200u
C9 GND VSS 2200u
C1 VDD GND 220n
C2 VDD GND 2200u
C3 VDD GND 2200u
C6 Net-_C17-Pad1_ /InL 1u
R3 Net-_C17-Pad1_ GNDA 22k
P2 GNDA /InL IN-L
R1 /OutL Net-_R1-Pad2_ 22k
R2 Net-_C5-Pad1_ Net-_R1-Pad2_ 680
C5 Net-_C5-Pad1_ GNDA 22u/25V
C4 Net-_C4-Pad1_ /OutL 22u/63V
P1 Net-_L1-Pad2_ GND OUT-L
P3 GND GND VDD VSS POWER
U2 GNDA Net-_R8-Pad2_ Net-_C16-Pad1_ GNDA Net-_C14-Pad1_ VDD VSS xStby xMute VDD /OutR VSS TDA7294V
C16 Net-_C16-Pad1_ /InR 1u
R10 Net-_C16-Pad1_ GNDA 22k
P6 GNDA /InR IN-R
R8 /OutR Net-_R8-Pad2_ 22k
R9 Net-_C15-Pad1_ Net-_R8-Pad2_ 680
C15 Net-_C15-Pad1_ GNDA 22u/25V
C14 Net-_C14-Pad1_ /OutR 22u/63V
P5 Net-_L2-Pad2_ GND OUT-R
P4 GNDA Net-_P4-Pad2_ MUTE
C10 xMute GNDA 10u
C11 xStby GNDA 10u
R15 Net-_D1-Pad1_ xMute 22k
R14 Net-_D1-Pad1_ xStby 10k
D1 Net-_D1-Pad1_ xMute 1N4148
R6 VDD Net-_Q1-Pad3_ 100k
R4 VDD Net-_P4-Pad2_ 47k
R5 Net-_P4-Pad2_ GNDA 47k
Q1 Net-_P4-Pad2_ GNDA Net-_Q1-Pad3_ BC846
Q2 Net-_Q1-Pad3_ GNDA Net-_Q2-Pad3_ BC846
R11 Net-_Q3-Pad1_ Net-_Q2-Pad3_ 68k
R7 VDD Net-_Q3-Pad1_ 30k
Q3 Net-_Q3-Pad1_ VDD Net-_Q3-Pad3_ BC856
R12 Net-_Q3-Pad3_ Net-_D1-Pad1_ 20k
Q4 Net-_P4-Pad2_ GNDA Net-_D1-Pad1_ BC846
R13 Net-_D1-Pad1_ GNDA *
C12 VDD GND 220n
C13 GND VSS 220n
L1 /OutL Net-_L1-Pad2_ L
C17 Net-_C17-Pad1_ /InL 1u
C18 Net-_C16-Pad1_ /InR 1u
R16 GND GNDA 47
L2 /OutR Net-_L2-Pad2_ L
.end
