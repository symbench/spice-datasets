.title KiCad schematic
U1 NC_01 NC_02 NC_03 NRST VDD Button NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 Buzzer NC_10 GND VDD NC_11 NC_12 SWDIO SWCLK STM32F042F4Px
J1 Button Buzzer GND VDD SWDIO SWCLK NRST Conn_01x07_Female
.end
