.title KiCad schematic
U4 Net-_R3-Pad2_ Net-_R2-Pad1_ NC_01 NC_02 NC_03 NC_04 +5V GND Net-_C5-Pad2_ Net-_C6-Pad1_ NC_05 NC_06 NC_07 NC_08 1VpO GATE_OUT NC_09 NC_10 NC_11 +5V NC_12 GND NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 ATmega328-PU
J1 NC_19 Net-_J1-Pad2_ NC_20 Net-_J1-Pad4_ NC_21 DIN-5
R1 Net-_R1-Pad1_ Net-_J1-Pad2_ 220
U3 Net-_R1-Pad1_ Net-_J1-Pad4_ NC_22 GND Net-_R2-Pad1_ NC_23 4N35
Y1 Net-_C5-Pad2_ Net-_C6-Pad1_ 16 MHz Crystal
C6 Net-_C6-Pad1_ GND 22pF
C5 GND Net-_C5-Pad2_ 22pF
R3 +5V Net-_R3-Pad2_ 10K
J5 Net-_D2-Pad1_ Net-_D2-Pad1_ GND GND GND GND GND GND Net-_D1-Pad2_ Net-_D1-Pad2_ Conn_01x10
D1 +12V Net-_D1-Pad2_ 1N4148
D2 Net-_D2-Pad1_ -12V 1N4148
U2 +12V GND +5V LM7805_TO220
R2 Net-_R2-Pad1_ +5V 1k
C1 +12V GND 10uF
C4 +5V GND 10uF
U1 Net-_R8-Pad1_ Net-_R8-Pad1_ Net-_C10-Pad2_ -12V GATE_OUT Net-_R9-Pad1_ Net-_R9-Pad1_ +12V TL072
C2 GND +12V 0.1uF
C7 +12V GND 10uF
C8 GND -12V 10uF
C3 -12V GND 0.1uF
R4 1VpO Net-_C10-Pad2_ 5.1k
C10 GND Net-_C10-Pad2_ 0.47uF
J4 GND Net-_J4-PadT_ NC_24 CV Note
J3 GND Net-_J3-PadT_ NC_25 Gate Out
D3 Net-_D3-Pad1_ Net-_D3-Pad2_ LED
Q1 GND Net-_Q1-Pad2_ Net-_D3-Pad1_ 2N3904
R7 +5V Net-_D3-Pad2_ 1K
R6 GATE_OUT Net-_Q1-Pad2_ 1K
C9 GND Net-_C10-Pad2_ 0.47uF
R5 GND GATE_OUT 1M
R9 Net-_R9-Pad1_ Net-_J3-PadT_ 1K
R8 Net-_R8-Pad1_ Net-_J4-PadT_ 1K
.end
