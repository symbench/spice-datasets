.title KiCad schematic
BackConnector1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 NC_43 NC_44 NC_45 NC_46 NC_47 NC_48 NC_49 NC_50 Conn_02x25_Odd_Even
Omnetics1 NC_51 NC_52 NC_53 NC_54 NC_55 NC_56 NC_57 NC_58 NC_59 NC_60 NC_61 NC_62 NC_63 NC_64 NC_65 NC_66 NC_67 NC_68 NC_69 NC_70 NC_71 NC_72 NC_73 NC_74 NC_75 NC_76 NC_77 NC_78 NC_79 NC_80 NC_81 NC_82 NC_83 NC_84 NC_85 NC_86 Conn_02x18_Odd_Even
.end
