.title KiCad schematic
U3 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 GND NC_12 NC_13 NC_14 NC_15 NC_16 Net-_U2-Pad14_ NC_17 Z80_~RD NC_18 NC_19 NC_20 VCC 6116
U1 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 GND NC_34 NC_35 NC_36 NC_37 NC_38 Net-_U1-Pad20_ NC_39 Z80_~RD NC_40 NC_41 NC_42 NC_43 VCC VCC Atmel 28C64
U2 NC_44 GND GND GND NC_45 NC_46 NC_47 GND NC_48 NC_49 NC_50 NC_51 NC_52 Net-_U2-Pad14_ Net-_U1-Pad20_ VCC 74HCT138
.end
