.title KiCad schematic
IC1 Net-_IC1-Pad1_ NC_01 NC_02 NC_03 NC_04 NC_05 Net-_IC1-Pad1_ LDL212PUR
.end
