.title KiCad schematic
U1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 ATTINY85-20PU
U2 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 ATTINY85-20SU
U3 NC_17 NC_18 NC_19 NC_20 NC_21 4011
.end
