.title KiCad schematic
U3 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 Terminus_Technology_FE2.1
.end
