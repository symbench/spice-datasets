.title KiCad schematic
C1 Net-_C1-Pad1_ V_out1 4.7uF
C2 Net-_C2-Pad1_ V_out1 2.2uF
C3 Net-_C3-Pad1_ V_out1 10uF
C4 Net-_C4-Pad1_ V_out1 4.7uF
C5 Net-_C5-Pad1_ V_out1 1uF
C6 Net-_C6-Pad1_ V_out1 330uF
C7 Net-_C7-Pad1_ V_out1 0.22uF
C8 Net-_C8-Pad1_ V_out1 10uF
R2 Net-_J13-Pad2_ V_out2 3.3k
R3 Net-_J14-Pad2_ V_out2 10k
R4 Net-_J15-Pad2_ V_out2 59k
R5 Net-_J16-Pad2_ V_out2 1k
R6 Net-_J17-Pad2_ V_out2 10k
R7 Net-_J18-Pad2_ V_out2 20k
R8 Net-_J19-Pad2_ V_out2 100k
R9 Net-_J20-Pad2_ V_out2 330
C10 Net-_C10-Pad1_ V_out1 10uF
C12 V_out2 GND 10uF
C9 Net-_C9-Pad1_ V_out1 0.22uF
R1 V_out1 GND 10k
C11 Net-_C11-Pad1_ V_out1 10uF
J1 V_in Net-_C1-Pad1_ Conn_01x02
J21 V_out2 GND Conn_01x02
J12 V_out1 GND Conn_01x02
J2 V_in Net-_C2-Pad1_ Conn_01x02
J3 V_in Net-_C3-Pad1_ Conn_01x02
J4 V_in Net-_C4-Pad1_ Conn_01x02
J5 V_in Net-_C5-Pad1_ Conn_01x02
J6 V_in Net-_C6-Pad1_ Conn_01x02
J7 V_in Net-_C7-Pad1_ Conn_01x02
J8 V_in Net-_C8-Pad1_ Conn_01x02
J9 V_in Net-_C9-Pad1_ Conn_01x02
J10 V_in Net-_C10-Pad1_ Conn_01x02
J11 V_in Net-_C11-Pad1_ Conn_01x02
J13 V_in Net-_J13-Pad2_ Conn_01x02
J14 V_in Net-_J14-Pad2_ Conn_01x02
J15 V_in Net-_J15-Pad2_ Conn_01x02
J16 V_in Net-_J16-Pad2_ Conn_01x02
J17 V_in Net-_J17-Pad2_ Conn_01x02
J18 V_in Net-_J18-Pad2_ Conn_01x02
J19 V_in Net-_J19-Pad2_ Conn_01x02
J20 V_in Net-_J20-Pad2_ Conn_01x02
J0 GND V_in Conn_01x02
.end
