.title KiCad schematic
J55 Net-_J54-Pad4_ Net-_J54-Pad3_ NC_01 Audio-Jack-3
J54 NC_02 NC_03 Net-_J54-Pad3_ Net-_J54-Pad4_ NC_04 NC_05 InConnector
J56 Net-_C172-Pad2_ NC_06 Net-_J56-Pad3_ Net-_J56-Pad4_ NC_07 Net-_C173-Pad1_ OutConnector
R302 Net-_R302-Pad1_ Net-_J56-Pad4_ R
R301 NC_08 Net-_J56-Pad4_ R
U33 Net-_J56-Pad4_ Net-_R302-Pad1_ Net-_C169-Pad1_ NC_09 Net-_C170-Pad1_ Net-_R303-Pad1_ Net-_J56-Pad3_ NC_10 ADA4807-2ARM
R303 Net-_R303-Pad1_ Net-_J56-Pad3_ R
R304 NC_11 Net-_J56-Pad3_ R
C172 NC_12 Net-_C172-Pad2_ C
C174 NC_13 Net-_C172-Pad2_ C
C173 Net-_C173-Pad1_ NC_14 C
C175 Net-_C173-Pad1_ NC_15 C
C169 Net-_C169-Pad1_ Net-_C169-Pad2_ C
C170 Net-_C170-Pad1_ Net-_C170-Pad2_ C
R299 Net-_C171-Pad2_ Net-_C169-Pad1_ R
R300 Net-_C170-Pad1_ Net-_C171-Pad2_ R
R297 NC_16 Net-_C171-Pad2_ 10k
R298 Net-_C171-Pad2_ NC_17 10k
C171 NC_18 Net-_C171-Pad2_ 10u
R295 Net-_J54-Pad3_ Net-_C169-Pad2_ 2k2
R296 Net-_J54-Pad4_ Net-_C170-Pad2_ 2k2
D7 NC_19 Net-_C169-Pad2_ D
D9 Net-_C169-Pad2_ NC_20 D
D8 NC_21 Net-_C170-Pad2_ D
D10 Net-_C170-Pad2_ NC_22 D
.end
