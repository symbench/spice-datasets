.title KiCad schematic
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 5.6u
R1 Net-_C1-Pad2_ 0 1k
V1 Net-_C1-Pad1_ 0 pulse(0 4 2m 1n 1n 2m 4m)
.end
