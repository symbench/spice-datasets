.title KiCad schematic
U1 GND SCL SDA Btn1 Btn3 Btn5 Btn7 Btn9 A1 A3 RST RX TX Btn2 Btn4 Btn6 Btn8 A0 A2 Vin CardEdge_2x10
J13 GND Btn1 CONN_01X02
J17 GND Btn1 CONN_01X02_FEMALE
J21 GND Btn1 CONN_01X02_MALE
J14 GND Btn2 CONN_01X02
J18 GND Btn2 CONN_01X02_FEMALE
J22 GND Btn2 CONN_01X02_MALE
J15 GND Btn3 CONN_01X02
J19 GND Btn3 CONN_01X02_FEMALE
J23 GND Btn3 CONN_01X02_MALE
J16 GND Btn4 CONN_01X02
J20 GND Btn4 CONN_01X02_FEMALE
J24 GND Btn4 CONN_01X02_MALE
J25 GND Btn5 CONN_01X02
J30 GND Btn5 CONN_01X02_FEMALE
J35 GND Btn5 CONN_01X02_MALE
J1 GND Vin CONN_01X02
J4 GND Vin CONN_01X02_FEMALE
J9 GND Vin CONN_01X02_MALE
J2 GND Vin CONN_01X02
J6 GND Vin CONN_01X02_FEMALE
J10 GND Vin CONN_01X02_MALE
J3 RX TX CONN_01X02
J7 RX TX CONN_01X02_FEMALE
J11 RX TX CONN_01X02_MALE
J5 SCL SDA CONN_01X02
J8 SCL SDA CONN_01X02_FEMALE
J12 SCL SDA CONN_01X02_MALE
J40 GND A0 Vin CONN_01X03
J48 GND A0 Vin CONN_01X03_MALE
J41 GND A1 Vin CONN_01X03
J49 GND A1 Vin CONN_01X03_MALE
J42 GND A2 Vin CONN_01X03
J50 GND A2 Vin CONN_01X03_MALE
J43 GND A3 Vin CONN_01X03
J51 GND A3 Vin CONN_01X03_MALE
U2 GND Btn6 SaB-Jmp
U3 GND Btn7 SaB-Jmp
U4 GND Btn8 SaB-Jmp
U5 GND Btn9 SaB-Jmp
J26 GND RST CONN_01X02
J27 GND RST CONN_01X02_FEMALE
J28 GND RST CONN_01X02_MALE
.end
