.title KiCad schematic
IC2 GND Net-_IC2-Pad2_ NC_01 Net-_IC2-Pad4_ VBAT BTS500601TEAAUMA2
TP1 NC_02 TestPoint
J6 GND NC_03 NC_04 Conn_01x03
J10 Net-_J10-Pad1_ GND GND GND GND PCB.MMCX.F.ST.SMT.JACK.HT
J8 TES-GPS-FLAG VBAT Conn_01x02
R21 +5V Net-_R21-Pad2_ 523k
C34 Net-_C34-Pad1_ GND 430pF
C33 +5V GND 47uF
U8 VBAT VBAT GND +5V +5V Net-_R21-Pad2_ Net-_R19-Pad1_ Net-_C34-Pad1_ GND TPS82140
IC1 TES-EN +5V GND +3V3 Net-_IC1-Pad5_ GND MCP1826T-3302E_DC
J9 GND GND Net-_J10-Pad1_ U.FL-R-SMT_10_
J7 GND TES-EN TES-GPS-FLAG Conn_01x03
R23 GND Net-_IC2-Pad4_ 1k
C1 +3V3 GND 1uF
R22 NC_05 Net-_IC2-Pad4_ 10k
R20 NC_06 Net-_IC2-Pad2_ 10k
C32 VBAT GND 10uF
R19 Net-_R19-Pad1_ +5V 100k
R24 Net-_R21-Pad2_ GND 100k
R25 +3V3 Net-_IC1-Pad5_ 1k
TP3 NC_07 TestPoint
TP5 NC_08 TestPoint
TP7 NC_09 TestPoint
TP2 +3V3 TestPoint
TP4 +5V TestPoint
TP6 NC_10 TestPoint
TP8 NC_11 TestPoint
.end
