.title KiCad schematic
U1 NC_01 NC_02 NC_03 NC_04 NC_05 /TEST_THING NC_06 LM741
P1 /TEST_THING CONN_01X01
.end
