.title KiCad schematic
U2 GND GND NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 GND NC_14 NC_15 NC_16 NC_17 JTAG_TCK NC_18 SOP2 SOP1 NC_19 NC_20 GND GND NC_21 GND Net-_U1-Pad1_ GND NC_22 SOP0 CC_nRESET Net-_R8-Pad1_ +3V3 GND Net-_R9-Pad1_ +3V3 NC_23 NC_24 GND STATUS_LED_1 NC_25 NC_26 NC_27 STATUS_LED_2 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 GND GND GND GND GND GND GND GND GND CC3220MODSFMOB
U1 Net-_U1-Pad1_ GND Net-_J4-Pad1_ GND DEA202450BT-1294C1-H
J4 Net-_J4-Pad1_ GND WIFI SMA
R4 SOP0 GND 100k
R5 SOP1 GND 100k
R7 SOP2 GND 100k
R3 JTAG_TCK GND 100k
R6 +3V3 CC_nRESET 10k
C3 CC_nRESET GND 0.1uF
R8 Net-_R8-Pad1_ +3V3 DNP
C1 +3V3 GND 100uF
C2 +3V3 GND 100uF
C4 +3V3 GND 0.1uF
C5 +3V3 GND 0.1uF
C6 +3V3 GND 0.1uF
R9 Net-_R9-Pad1_ +3V3 DNP
R2 Net-_Q2-Pad3_ Net-_D6-Pad1_ 270
D6 Net-_D6-Pad1_ +3V3 LED
Q2 STATUS_LED_1 GND Net-_Q2-Pad3_ BSS138
R13 GND STATUS_LED_1 100k
R1 Net-_Q1-Pad3_ Net-_D5-Pad1_ 270
D5 Net-_D5-Pad1_ +3V3 LED
Q1 STATUS_LED_2 GND Net-_Q1-Pad3_ BSS138
R10 GND STATUS_LED_2 100k
.end
