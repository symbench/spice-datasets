.title KiCad schematic
J1 GND VCC IO13=RX IO14=TX Conn_01x04_Female
C1 VCC GND 10uF
C2 +3V3 GND 10uF
AE1 Net-_AE1-Pad1_ Net-_AE1-Pad2_ Antenna_Dipole
SW1 GND IO0=SW1 SW_Push
C3 +3V3 GND 100uF
U2 GND IO4=MISO IO12=MOSI IO27=SCK IO26=NSS IO25=RESET IO34=DIO5 GND Net-_AE1-Pad1_ Net-_AE1-Pad2_ IO21=DIO3 IO19=DIO4 +3V3 IO5=DIO0 IO17=DIO1 IO16=DIO2 RFM98W-433S2
U1 GND +3V3 +3V3 NC_01 NC_02 IO34=DIO5 NC_03 NC_04 NC_05 IO25=RESET IO26=NSS IO27=SCK IO14=TX IO12=MOSI GND IO13=RX NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 IO15=A NC_12 IO0=SW1 IO4=MISO IO16=DIO2 IO17=DIO1 IO5=DIO0 IO18=LED_RGB IO19=DIO4 NC_13 IO21=DIO3 RX0 TX0 NC_14 NC_15 GND GND ESP32-WROOM
U3 GND +3V3 VCC AMS1117-3.3
J2 GND +3V3 TX0 RX0 Conn_01x04_Female
J3 IO15=A Conn_01x01_Female
D1 /LED_VDD NC_16 GND IO18=LED_RGB WS2812B
R1 +3V3 /LED_VDD 75
.end
