.title KiCad schematic
U1 Net-_C9-Pad1_ Net-_C10-Pad1_ NC_01 /AREF NC_02 Net-_C7-Pad1_ NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 +3V3 Net-_U1-Pad18_ NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 Net-_U1-Pad18_ +3V3 NC_29 NC_30 NC_31 /~RESET_SAMD NC_32 Net-_U1-Pad18_ Net-_C6-Pad1_ NC_33 /SWCLK /SWDIO NC_34 NC_35 ATSAMD21G18A-AUT-MCU_Microchip_SAMD_Redone
C1 +3V3 GND 0.1uF
C2 +3V3 GND 10uF
C3 /AREF GND 1uF
C5 +3V3 GND 0.1uF
C4 +3V3 GND 10uF
C6 Net-_C6-Pad1_ GND 1uF
C7 Net-_C7-Pad1_ GND 10uF
C8 Net-_C7-Pad1_ GND 0.1uF
L1 +3V3 Net-_C7-Pad1_ 10uH
Y1 Net-_C9-Pad1_ Net-_C10-Pad1_ 32768Hz
C9 Net-_C9-Pad1_ GND 10pF
C10 Net-_C10-Pad1_ GND 10pF
TP1 /SWCLK TestPoint
TP2 /SWDIO TestPoint
SW1 /~RESET_SAMD GND SW_SPST
.end
