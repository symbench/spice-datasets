.title KiCad schematic
C5 Net-_C5-Pad1_ GND 2.2u
C3 Net-_C3-Pad1_ GND 6p
C4 Net-_C4-Pad1_ GND 6p
Y1 Net-_C4-Pad1_ Net-_C3-Pad1_ 8M
C8 +3V3 GND 0.1u
C10 +3V3 GND 0.1u
C12 +3V3 GND 0.1u
C13 +3V3 GND 0.1u
C14 +3V3 GND 0.1u
C15 +3V3 GND 4.7u
C6 +3V3 GND 0.1u
C7 +3V3 GND 0.1u
C9 +3V3 GND 1u
C11 /NRST GND 0.1u
SW1 /NRST GND Reset
J3 +3V3 /SWCLK /SWDIO GND SWD
J2 +3V3 Net-_J2-Pad2_ GND Bootloader
U1 NC_01 NC_02 GND /D+ /D- +3V3 +3V3 Net-_R1-Pad1_ Net-_R2-Pad2_ NC_03 NC_04 GND NC_05 NC_06 /USART2_RTS /USART2_CTS /USART2_TX /USART2_RX NC_07 NC_08 GND CP2102N-A01-GQFN20
R2 +3V3 Net-_R2-Pad2_ 1k
C2 +3V3 GND 4.7u
C1 +3V3 GND 0.1u
R3 GND Net-_R1-Pad1_ 47.5k
R1 Net-_R1-Pad1_ +5V 22.k
J1 GND +5V Net-_J1-PadA5_ /D+ /D- NC_09 +5V GND GND +5V Net-_J1-PadB5_ /D+ /D- NC_10 +5V GND GND USB_C_Receptacle_USB2.0
D1 GND /D+ /D- +5V SP0503BAHT
R4 Net-_J1-PadB5_ GND 5.1k
R5 Net-_J1-PadA5_ GND 5.1k
U2 +3V3 NC_11 NC_12 NC_13 Net-_C3-Pad1_ Net-_C4-Pad1_ /NRST NC_14 NC_15 NC_16 NC_17 GND +3V3 /USART2_CTS /USART2_RTS /USART2_TX /USART2_RX GND +3V3 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 Net-_C5-Pad1_ GND +3V3 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 /SWDIO GND +3V3 /SWCLK NC_41 NC_42 NC_43 NC_44 NC_45 NC_46 NC_47 NC_48 NC_49 NC_50 Net-_J2-Pad2_ NC_51 NC_52 GND +3V3 STM32F413RHTx
.end
