.title KiCad schematic
U5 NC_01 NC_02 NC_03 Net-_U5-Pad4_ NC_04 NC_05 NC_06 Net-_U5-Pad4_ NC_07 TP4056
.end
