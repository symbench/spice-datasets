.title KiCad schematic
X2 NC_01 GND NC_02 NC_03 NC_04 NC_05 GND GND MAB6H
C1 5V0 GND 100nF
C3 GND 3V3_PWR6 100nF
.end
