.title KiCad schematic
JS1 JS1_1 JS1_2 JS1_3 JS1_4 JS1_5 JS1_6 JS1_7 GND JS1_9 Serial Port
R8 JS1_5 3V3_PWR6 47K
R6 JS1_4 3V3_PWR6 47K
R5 JS1_3 3V3_PWR6 47K
R3 JS1_2 3V3_PWR6 47K
R1 JS1_1 3V3_PWR6 47K
R2 JS1_6 3V3_PWR6 47K
R4 JS1_7 3V3_PWR6 47K
R7 JS1_9 3V3_PWR6 47K
JS2 JS2_1 JS2_2 JS2_3 JS2_4 JS2_5 JS2_6 JS2_7 GND JS2_9 Serial Port
R12 JS2_5 JOY_3V3 47K
R13 JS2_4 JOY_3V3 47K
R14 JS2_3 JOY_3V3 47K
R15 JS2_2 JOY_3V3 47K
R16 JS2_1 JOY_3V3 47K
R19 JS2_6 JOY_3V3 47K
R20 JS2_7 JOY_3V3 47K
R21 JS2_9 JOY_3V3 47K
.end
