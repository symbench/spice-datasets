.title KiCad schematic
U1 GND G11 PCM_CLK PCM_FS G17 G16 G15 Net-_J6-Pad2_ Net-_J6-Pad3_ MISO MOSI SCK CS PCM_DOUT PCM_DIN RST SDA SCL G19 G18 /E_RX+ /E_RX- /E_TX+ /E_TX- VCCQ FW_RST Net-_J5-Pad3_ Net-_J5-Pad2_ /U_D- /U_D+ +3V3 GND Omega2+
J3 +3V3 GND Conn_01x02
J5 GND Net-_J5-Pad2_ Net-_J5-Pad3_ UART0
J6 GND Net-_J6-Pad2_ Net-_J6-Pad3_ UART1
J7 VCCQ /E_TX- /E_TX+ /E_RX- /E_RX+ GND GND ETH
J4 +3V3 SDA SCL G17 GND I2C
J2 GND /U_D- /U_D+ +3V3 GND USB
J1 MOSI MISO SCK CS +3V3 GND PCM_CLK PCM_DIN PCM_DOUT PCM_FS GND +5V Conn_01x12
SW2 Net-_R1-Pad2_ FW_RST FW_RST
R1 +3V3 Net-_R1-Pad2_ 1K
SW1 GND RST RST
J8 +3V3 G15 G16 G17 G11 G18 G19 GND Conn_01x08
.end
