.title KiCad schematic
C12 /V_DEVICE GND 4.7u
C10 VDD GND 4.7u
C9 VDD GND 100n
U1 /SCL /INTB /PORT /A+ /A- VDD /B- /B+ /ID /VCONN /CC1 /CC2 /ENB /B1+ /B1- /A1+ /A1- /B2- /B2+ /A2- /A2+ /ADDR Net-_R2-Pad1_ /SDA GND PI5USB30213A
C8 /A2+ /TX2+ 100n
C7 /A2- /TX2- 100n
C6 /B2+ /RX2+ 100n
C5 /B2- /RX2- 100n
C4 /A1+ /TX1+ 100n
C3 /A1- /TX1- 100n
C2 /B1+ /RX1+ 100n
R1 VDD VBUS 0R
R2 Net-_R2-Pad1_ VBUS 910K
C1 /B1- /RX1- 100n
J6 /V_DEVICE /D- /D+ GND /SSRX- /SSRX+ GND /SSTX- /SSTX+ GND USB3_A
J1 GND /TX1+ /TX1- VBUS /CC1 /D+ /D- Net-_J1-PadA8_ VBUS /RX2- /RX2+ GND GND /TX2+ /TX2- VBUS /CC2 /D+ /D- Net-_J1-PadB8_ VBUS /RX1- /RX1+ GND GND USB_C_Receptacle
R5 /SSTX- /A- 0R
R6 /SSTX+ /A+ 0R
C13 /SSRX- /B- 100n
C14 /SSRX+ /B+ 100n
R12 VDD Net-_J5-Pad17_ 1K
R13 VDD Net-_J5-Pad15_ 4K7
R14 GND Net-_J5-Pad11_ 4K7
R15 VDD Net-_J5-Pad9_ 4K7
R16 GND Net-_J5-Pad5_ 4K7
J2 /TX1- /TX1+ GND /RX1- /RX1+ /RX1+ /RX1- GND /TX1+ /TX1- PUSB3FR4Z
J4 /TX2+ /TX2- GND /RX2+ /RX2- /RX2- /RX2+ GND /TX2- /TX2+ PUSB3FR4Z
J8 /ID /SCL /SDA /INTB Conn_IO
R8 /SDA Net-_J5-Pad29_ 2.2K
R9 /SCL Net-_J5-Pad27_ 2.2K
R10 /ID Net-_J5-Pad25_ 2.2K
R7 /INTB Net-_J5-Pad31_ 2.2K
SBU1 Net-_J1-PadA8_ TestPoint
SBU2 Net-_J1-PadB8_ TestPoint
J5 /CC1 /CC1 /CC2 /CC2 Net-_J5-Pad5_ /PORT NC_01 /PORT Net-_J5-Pad9_ /PORT Net-_J5-Pad11_ /ADDR NC_02 /ADDR Net-_J5-Pad15_ /ADDR Net-_J5-Pad17_ /ENB /V_DEVICE /VCONN /V_DEVICE /VCONN /V_DEVICE VDD Net-_J5-Pad25_ VDD Net-_J5-Pad27_ VDD Net-_J5-Pad29_ VDD Net-_J5-Pad31_ VDD VDD VDD GND GND 02x18
.end
