.title KiCad schematic
J1 /A0 /A1 /A2 /A3 /A4 /A5 /A6 /A7 /A8 /A9 /A10 /A11 /A12 /A13 /A14 /A15 /A16 /A17 /A18 /A19-IO15 /~CE1 /CE2 Conn_01x22_Male
J2 GND +3V3 ~BLE ~BHE ~BYTE ~OE ~WE /IO14 /IO13 /IO12 /IO11 /IO10 /IO9 /IO8 /IO7 /IO6 /IO5 /IO4 /IO3 /IO2 /I01 /IO0 Conn_01x22_Male
C1 GND +3V3 0.1uF
U1 /A15 /A14 /A13 /A12 /A11 /A10 /A9 /A8 NC_01 NC_02 ~WE /CE2 NC_03 ~BHE ~BLE /A18 /A17 /A7 /A6 /A5 /A4 /A3 /A2 /A1 /A0 /~CE1 GND ~OE /IO0 /IO8 /I01 /IO9 /IO2 /IO10 /IO3 /IO11 +3V3 /IO4 /IO12 /IO5 /IO13 /IO6 /IO14 /IO7 /A19-IO15 GND ~BYTE /A16 CY62157
.end
