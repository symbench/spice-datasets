.title KiCad schematic
SW1 ROW3 Net-_D1-Pad1_ 7
D1 Net-_D1-Pad1_ COL0 DIODE
SW2 ROW3 Net-_D2-Pad1_ 8
D2 Net-_D2-Pad1_ COL1 DIODE
SW3 ROW3 Net-_D3-Pad1_ 9
D3 Net-_D3-Pad1_ COL2 DIODE
SW5 ROW2 Net-_D5-Pad1_ 4
D5 Net-_D5-Pad1_ COL0 DIODE
SW6 ROW2 Net-_D6-Pad1_ 5
D6 Net-_D6-Pad1_ COL1 DIODE
SW7 ROW2 Net-_D7-Pad1_ 6
D7 Net-_D7-Pad1_ COL2 DIODE
SW9 ROW1 Net-_D9-Pad1_ 1
D9 Net-_D9-Pad1_ COL0 DIODE
SW13 ROW0 Net-_D13-Pad1_ 0
D13 Net-_D13-Pad1_ COL0 DIODE
SW10 ROW1 Net-_D10-Pad1_ 2
D10 Net-_D10-Pad1_ COL1 DIODE
SW14 ROW0 Net-_D14-Pad1_ .
D14 Net-_D14-Pad1_ COL1 DIODE
SW11 ROW1 Net-_D11-Pad1_ 3
D11 Net-_D11-Pad1_ COL2 DIODE
SW15 ROW0 Net-_D15-Pad1_ /
D15 Net-_D15-Pad1_ COL2 DIODE
SW4 ROW3 Net-_D4-Pad1_ -
D4 Net-_D4-Pad1_ COL3 DIODE
SW8 ROW2 Net-_D8-Pad1_ *
D8 Net-_D8-Pad1_ COL3 DIODE
SW12 ROW1 Net-_D12-Pad1_ +
D12 Net-_D12-Pad1_ COL3 DIODE
SW16 ROW0 Net-_D16-Pad1_ Enter
D16 Net-_D16-Pad1_ COL3 DIODE
U1 GND NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 ROW4 COL0 COL1 COL2 COL3 ROW0 ROW1 ROW2 ROW3 NC_18 NC_19 NC_20 NC_21 Teensy2.0
SW17 ROW4 Net-_D17-Pad1_ Blank1
D17 Net-_D17-Pad1_ COL0 DIODE
SW18 ROW4 Net-_D18-Pad1_ Blank2
D18 Net-_D18-Pad1_ COL1 DIODE
H1 GND MountingHole_Pad
H8 GND MountingHole_Pad
H7 GND MountingHole_Pad
H6 GND MountingHole_Pad
H5 GND MountingHole_Pad
H4 GND MountingHole_Pad
H3 GND MountingHole_Pad
H2 GND MountingHole_Pad
.end
