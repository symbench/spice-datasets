.title KiCad schematic
U1 /RA5 NC_01 /MCLR /RC5 /RC4 /RC3 /RC2 /RC1 /RC0 NC_02 /ICSPCLK /ICSPDAT GND NC_03 NC_04 +BATT GND PIC16F1503_QFN
D4 /RC0 Net-_D4-PadC_ LED_0603
D3 /RC0 Net-_D3-PadC_ LED_0603
D2 /RC0 Net-_D2-PadC_ LED_0603
D7 /RC1 Net-_D7-PadC_ LED_0603
D6 /RC1 Net-_D6-PadC_ LED_0603
D5 /RC1 Net-_D5-PadC_ LED_0603
D10 /RC2 Net-_D10-PadC_ LED_0603
D9 /RC2 Net-_D9-PadC_ LED_0603
D8 /RC2 Net-_D8-PadC_ LED_0603
R5 Net-_D4-PadC_ /RC5 RES_0603
R4 Net-_D3-PadC_ /RC4 RES_0603
R3 Net-_D2-PadC_ /RC3 RES_0603
R8 Net-_D7-PadC_ /RC5 RES_0603
R7 Net-_D6-PadC_ /RC4 RES_0603
R6 Net-_D5-PadC_ /RC3 RES_0603
R11 Net-_D10-PadC_ /RC5 RES_0603
R10 Net-_D9-PadC_ /RC4 RES_0603
R9 Net-_D8-PadC_ /RC3 RES_0603
C2 +BATT GND CAP_0603
J1 /MCLR Net-_J1-Pad2_ GND /ICSPDAT /ICSPCLK NC_05 HEADER_1X6
R1 Net-_C1-Pad1_ +BATT RES_0603
C1 Net-_C1-Pad1_ GND CAP_0603
D1 Net-_C1-Pad1_ /MCLR Schottky_SMA
R2 +BATT Net-_J1-Pad2_ RES_0603
SW1 GND Net-_R12-Pad1_ SWITCH_MOMENTARY
R12 Net-_R12-Pad1_ /RA5 RES_0603
.end
