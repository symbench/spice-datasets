.title KiCad schematic
J2 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 Digital pins
J4 NC_10 NC_11 NC_12 NC_13 I2C
J3 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 ICSP
J1 NC_20 NC_21 NC_22 NC_23 Serial
.end
