.title KiCad schematic
U201 NC_01 NC_02 /EMMC_DAT7 /EMMC_DAT6 /EMMC_DAT2 /~EMMC_RST NC_03 /EMMC_DAT5 /EMMC_DAT1 NC_04 /EMMC_DAT4 Net-_R403-Pad1_ NC_05 /EMMC_DAT3 /EMMC_DAT0 Net-_R402-Pad1_ NC_06 PP_NAND_IO MCIMX6Y2DVM
U401 Net-_C407-Pad1_ PP_NAND_FLASH PP_NAND_FLASH PP_NAND_FLASH PP_NAND_FLASH PP_NAND_FLASH PP_NAND_FLASH PP_NAND_FLASH PP_NAND_FLASH COM COM COM COM COM COM COM COM COM PP_NAND_IO PP_NAND_IO COM /EMMC_DAT0 /EMMC_DAT2 /EMMC_DAT5 /EMMC_DAT7 PP_NAND_IO COM PP_NAND_IO PP_NAND_IO COM PP_NAND_IO COM /~EMMC_RST COM /EMMC_DAT1 /EMMC_DAT3 /EMMC_DAT4 /EMMC_DAT6 COM PP_NAND_IO /EMMC_CMD /EMMC_CLK PP_NAND_IO COM MTFC8GACAANA-4M
C402 PP_NAND_IO COM 0.22u
C401 PP_NAND_IO COM 10u
C404 PP_NAND_FLASH COM 0.22u
C403 PP_NAND_FLASH COM 10u
C408 Net-_C407-Pad1_ COM 0.22u
C407 Net-_C407-Pad1_ COM 10u
R402 Net-_R402-Pad1_ /EMMC_CLK 22
C406 PP_NAND_IO COM 0.22u
C405 PP_NAND_IO COM 10u
R403 Net-_R403-Pad1_ /EMMC_CMD 22
R401 /~EMMC_RST COM 10k
.end
