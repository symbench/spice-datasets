.title KiCad schematic
A1 BT_RX BT_TX NC_01 GND NEO PWM_DER I2C_SDA I2C_SCL PWM_IZQ D7 D8 D9 D10 D11 LINEA_SEL D13 NC_02 NC_03 BAT A1 LINEA_1 LINEA_2 LINEA_3 DIST_DCHA DIST_FRONT DIST_IZQ +5V NC_04 GND VCC Arduino_Nano_v3.x
J7 VBAT NC_05 GND Conn_01x03
J8 Net-_J8-Pad1_ GND Conn_01x02
J9 VBAT Net-_J8-Pad1_ Conn_01x02
R3 +5V Net-_D2-Pad2_ R
R4 +5V Net-_D3-Pad2_ R
D2 LED_R Net-_D2-Pad2_ LED
D3 LED_G Net-_D3-Pad2_ LED
R5 +5V B1 R
R6 +5V B2 R
SW1 B1 GND SW_Push
SW2 B2 GND SW_Push
U2 GND GND GND LED_G LED_R DIR_IZQ_1 DIR_IZQ_2 GND DIR_DER_1 DIR_DER_2 B1 B2 NC_06 I2C_SCL I2C_SDA +5V PCF8574
R8 +5V I2C_SDA R
R7 +5V I2C_SCL R
J6 D7 D8 D9 Conn_01x03
J5 D10 D11 D13 Conn_01x03
J10 A1 +5V +5V Conn_01x03
J11 GND GND GND Conn_01x03
J12 NC_07 +5V GND Net-_D4-Pad1_ BT_RX NC_08 Conn_01x06
D4 Net-_D4-Pad1_ BT_TX D
SW3 NC_09 VBAT VDD NC_10 +5V STBY_MOT SW_DPDT_x2
JP1 VDD VCC Jumper_NO_Small
D5 Net-_D5-Pad1_ GND +5V NEO NeoPixel_THT
D6 NC_11 GND +5V Net-_D5-Pad1_ NeoPixel_THT
C1 GND +5V C
C2 GND +5V C
J4 PWM_IZQ DIR_IZQ_2 DIR_IZQ_1 STBY_MOT DIR_DER_1 DIR_DER_2 PWM_DER GND Conn_01x08
J1 VBAT +5V GND M_IXQ_+ M_IXQ_- M_DER_- M_DER_+ GND Conn_01x08
J2 M_IXQ_- M_IXQ_+ Conn_01x02
J3 M_DER_- M_DER_+ Conn_01x02
R1 VDD BAT R_Small
R2 BAT GND R_Small
D1 +5V BAT D_Small
J13 +5V GND LINEA_1 LINEA_2 LINEA_3 LINEA_SEL Conn_01x06
J14 DIST_IZQ GND +5V Conn_01x03
J15 DIST_FRONT GND +5V Conn_01x03
J16 DIST_DCHA GND +5V Conn_01x03
U1 VDD GND +5V GND DC-DC_BuckModule
.end
