.title KiCad schematic
U4 +9V GND +5V L7805
U2 +5V /ESP32_RX_5V /ESP32_TX GND /PIC32_RX /PIC32_~RX /PIC32_~TX /PIC32_TX SN75179BD
R1 /ESP32_RX_3V3 /ESP32_RX_5V 1K
D2 +3V3 /ESP32_RX_3V3 1N4148
D5 Net-_D5-Pad1_ Net-_D5-Pad2_ LED
D3 Net-_D3-Pad1_ Net-_D3-Pad2_ LED
R2 Net-_D3-Pad1_ GND 220
R4 Net-_D5-Pad1_ GND 220
U3 +3V3 NC_01 NC_02 NC_03 /GPIO0 /GPIO15 Net-_D3-Pad2_ Net-_D5-Pad2_ /ESP32_RX_3V3 /ESP32_TX NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 +9V GND NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 DoitESP32-DevKit-V1
U1 Net-_C1-Pad1_ GND +9V L7809
C2 +9V GND 0.1uF 16V
C3 +5V GND 0.1uF 16V
C1 Net-_C1-Pad1_ GND 0.33uF 50v
J1 +3V3 +5V +9V GND /GPIO0 /GPIO15 Conn_01x06_Female
D1 Net-_C1-Pad1_ /15V_UnProtected B120-E3
D4 GND Net-_D4-Pad2_ LED
R3 +5V Net-_D4-Pad2_ 470
J2 GND NC_28 NC_29 NC_30 /15V_UnProtected GND /PIC32_RX /PIC32_~RX /PIC32_~TX /PIC32_TX DB9_Female_MountingHoles
.end
