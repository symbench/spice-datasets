.title KiCad schematic
J1 Net-_J1-Pad1_ Net-_J1-Pad1_ Net-_J1-Pad1_ Net-_J1-Pad1_ Net-_J1-Pad1_ Net-_J1-Pad1_ Net-_J1-Pad1_ Conn_01x07_Female
.end
