.title KiCad schematic
J1 5V GND 5V GND 5V GND 5V GND 5V GND 5V GND 5V GND NC_01 GND NC_02 NC_03 NC_04 NC_05 2X10-2MMSMD
.end
