.title KiCad schematic
H1 GND MountingHole_Pad
H2 GND MountingHole_Pad
U2 SCL SDA NC_01 3.3V GND NRST CH1_DATA CH2_DATA CH3_DATA NC_02 CH3_RX_EN CH3_TX_EN CH2_RX_EN CH2_TX_EN Net-_U1-Pad4_ CH1_RX_EN CH1_TX_EN SWDIO SWCLK COM_DATA STM32G030F6P6
R3 3.3V NRST R_US
SW1 GND NRST SW_Push
R1 3.3V SCL R_US
R2 3.3V SDA R_US
U1 5V GND LED_OUT Net-_U1-Pad4_ GND 3.3V SN74LVC1T45DBVR
J1 3.3V GND NRST SWDIO SWCLK Conn_01x05
J3 PRI_HI PRI_LO Conn_01x02
J4 PRI_HI PRI_LO Conn_01x02
J2 PRI_HI PRI_LO Conn_01x02
J5 CH1_DATA CH2_DATA CH3_DATA Conn_01x03
J6 LED_OUT GND 5V Conn_01x03
U3 CH1_TX_EN COM_DATA GND CH1_DATA 3.3V 74LVC1G125
U4 CH1_RX_EN CH1_DATA GND COM_DATA 3.3V 74LVC1G125
U5 CH2_TX_EN COM_DATA GND CH2_DATA 3.3V 74LVC1G125
U6 CH2_RX_EN CH2_DATA GND COM_DATA 3.3V 74LVC1G125
U7 CH3_TX_EN COM_DATA GND CH3_DATA 3.3V 74LVC1G125
U8 CH3_RX_EN CH3_DATA GND COM_DATA 3.3V 74LVC1G125
U9 3.3V 3.3V 3.3V GND SDA SCL GND 3.3V MB85RC256
C1 +VDC GND 10u
C2 +VDC GND 1u
C3 +VDC GND 0.1u
U11 5V GND 5V NC_03 3.3V AP2112K-3.3
C4 5V GND 0.1u
C5 3.3V GND 1u
U10 GND 5V +VDC LM1085-5.0
C6 3.3V GND 4.7u
CR1 +VDC GND PRI_LO PRI_HI DF01S
.end
