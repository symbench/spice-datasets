.title KiCad schematic
J1 GND /VCC Net-_J1-Pad3_ Net-_J1-Pad4_ Net-_J1-Pad5_ Net-_J1-Pad6_ Net-_J1-Pad7_ Net-_J1-Pad8_ Conn_01x08_Male
R2 Net-_J1-Pad3_ Net-_R2-Pad2_ 1K
R1 Net-_J1-Pad3_ /VCC 100
SW1 Net-_R2-Pad2_ GND up
R4 Net-_J1-Pad4_ Net-_R4-Pad2_ 1K
R3 Net-_J1-Pad4_ /VCC 100
SW2 Net-_R4-Pad2_ GND down
R6 Net-_J1-Pad5_ Net-_R6-Pad2_ 1K
R5 Net-_J1-Pad5_ /VCC 100
SW3 Net-_R6-Pad2_ GND right
R8 Net-_J1-Pad6_ Net-_R8-Pad2_ 1K
R7 Net-_J1-Pad6_ /VCC 100
SW4 Net-_R8-Pad2_ GND left
R10 Net-_J1-Pad7_ Net-_R10-Pad2_ 1K
R9 Net-_J1-Pad7_ /VCC 100
SW5 Net-_R10-Pad2_ GND confirm
R12 Net-_J1-Pad8_ Net-_R12-Pad2_ 1K
R11 Net-_J1-Pad8_ /VCC 100
SW6 Net-_R12-Pad2_ GND return
.end
