.title KiCad schematic
U1 GLV- NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 SPAN02A-12
.end
