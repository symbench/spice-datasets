.title KiCad schematic
J1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 USB_B_Micro
.end
