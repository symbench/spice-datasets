.title KiCad schematic
U1 NC_01 NC_02 NC_03 NC_04 NC_05 Net-_R2-Pad2_ Net-_R1-Pad2_ NC_06 GND NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 GND NC_13 NC_14 NC_15 NC_16 GND LT3751
U2 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 ACPL-C87B-000E
Q1 NC_25 NC_26 NC_27 NTB35N15
D1 NC_28 NC_29 RFN5TF8S
C1 +24V GND C
C2 +24V GND C
C3 +24V GND C
T1 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 +24V +24V +24V +24V GA3460-BL
C5 +24V GND C_2.2uF
C6 NC_38 NC_39 C_10uF_450V
R2 VCC Net-_R2-Pad2_ R_100K
R1 VCC Net-_R1-Pad2_ R_100K
C4 +24V GND C
R3 NC_40 NC_41 R_0
.end
