.title KiCad schematic
U1 GND Net-_L1-Pad1_ /V_down_1/12VIN Net-_C4-Pad2_ NC_01 Net-_C3-Pad2_ TPS563200
J1 GND /V_down_1/12VIN Conn_01x02_Female
L1 Net-_L1-Pad1_ /USB_1/5VIN 4.7uH
C3 /USB_1/5VIN Net-_C3-Pad2_ 0.1uF
R1 /USB_1/5VIN Net-_C4-Pad2_ 54.9k
R2 Net-_C4-Pad2_ GND 10k
C4 /USB_1/5VIN Net-_C4-Pad2_ 0.1uF
C5 Net-_C4-Pad2_ GND 0.1uF
C2 /V_down_1/12VIN GND 10uF
C1 /V_down_1/12VIN GND C
J2 /USB_1/USB_1_SUPPLY Net-_J2-Pad2_ Net-_J2-Pad3_ GND GND USB_A
U3 Net-_J2-Pad3_ GND Net-_J3-Pad3_ Net-_J3-Pad2_ /USB_1/5VIN Net-_J2-Pad2_ TPS2513A
U2 GND /USB_1/5VIN /USB_1/5VIN /USB_1/~FAULT1 /USB_1/~FAULT2 /USB_1/~FAULT1 Net-_R5-Pad1_ /USB_1/USB_2_SUPPLY /USB_1/USB_1_SUPPLY /USB_1/~FAULT2 GND TPS2561A
J3 /USB_1/USB_2_SUPPLY Net-_J3-Pad2_ Net-_J3-Pad3_ GND GND USB_A
C10 /USB_1/USB_1_SUPPLY GND CP1
C9 /USB_1/USB_2_SUPPLY GND CP1
R5 Net-_R5-Pad1_ GND 25.5K
C6 /USB_1/5VIN GND C
R3 /USB_1/5VIN /USB_1/~FAULT1 R
R4 /USB_1/5VIN /USB_1/~FAULT2 R
C7 /USB_1/~FAULT1 GND 0.22uF
C8 /USB_1/~FAULT2 GND 0.22uF
.end
