.title KiCad schematic
J1 GND VCC IO13=RX IO14=TX Conn_01x04_Female
C1 VCC GND 10uF
C2 +3V3 GND 10uF
SW1 GND IO0=SW1 SW_Push
C3 +3V3 GND 100uF
U1 GND +3V3 +3V3 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 IO25=SCK IO26=MOSI IO27=MISO IO14=TX NC_07 GND IO13=RX NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 IO15=A NC_14 IO0=SW1 IO4=DIO3 IO16=DIO2 IO17=DIO1 IO5=BUSY IO18=NRESET IO19=TX_EN NC_15 IO21=NSS RX0 TX0 IO22=RX_EN IO23=RGBLED GND GND ESP32-WROOM
U3 GND +3V3 VCC AMS1117-3.3
J2 GND +3V3 TX0 RX0 Conn_01x04_Female
J3 IO15=A Conn_01x01_Female
D1 /LED_VDD NC_16 GND IO23=RGBLED WS2812B
R1 +3V3 /LED_VDD 75
U2 +3V3 GND IO27=MISO IO26=MOSI IO25=SCK IO21=NSS GND IO22=RX_EN IO19=TX_EN GND IO18=NRESET IO5=BUSY IO17=DIO1 IO16=DIO2 IO4=DIO3 GND E28-2G4M20S
.end
