.title KiCad schematic
U1 Net-_P2-Pad2_ Net-_P2-Pad2_ Net-_RV1-Pad2_ Net-_RV1-Pad1_ Net-_P2-Pad1_ Net-_P2-Pad2_ Net-_P2-Pad2_ Net-_P2-Pad1_ Net-_RV1-Pad1_ Net-_RV1-Pad2_ Net-_P3-Pad2_ Net-_P3-Pad2_ Recom
RV1 Net-_RV1-Pad1_ Net-_RV1-Pad2_ Net-_P2-Pad1_ POT
P1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 CONN_01X19
P2 Net-_P2-Pad1_ Net-_P2-Pad2_ BNC
P3 Net-_P2-Pad2_ Net-_P3-Pad2_ NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 CONN_01X19
.end
