.title KiCad schematic
Motor11 NC_01 Stepper_motor_14HM11-0404S
.end
