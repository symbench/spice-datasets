.title KiCad schematic
M1 NC_01 NC_02 NC_03 NC_04 NC_05 DC_Motor
.end
