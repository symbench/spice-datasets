.title KiCad schematic
R1 +3V3 Net-_R1-Pad2_ 10k
P3 /TX /RX GND CONN_01X03
P2 /SCLK /MOSI /MISO /CSO CONN_01X04
P1 /ADC /GPIO16 /GPIO14 /GPIO12 /GPIO13 /GPIO5 /GPIO4 /GPIO0 /GPIO2 /GPIO15 /GPIO9 /GPIO10 CONN_01X12
P4 +3V3 GND CONN_01X02
FLSH1 /GPIO0 GND SW_PUSH
RST1 Net-_R1-Pad2_ GND SW_PUSH
R2 GND /GPIO15 10k
R3 +3V3 /GPIO2 10k
R4 +3V3 /GPIO0 10k
U1 Net-_R1-Pad2_ /ADC +3V3 /GPIO16 /GPIO14 /GPIO12 /GPIO13 +3V3 /CSO /MISO /GPIO9 /GPIO10 /MOSI /SCLK GND /GPIO15 /GPIO2 /GPIO0 /GPIO4 /GPIO5 /RX /TX ESP-12F
.end
