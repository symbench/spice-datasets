.title KiCad schematic
Q1 Net-_D1-Pad2_ NC_01 +24V Q_PMOS_GDS
D1 +24V Net-_D1-Pad2_ D_Zener
R1 Net-_D1-Pad2_ GND R
U1 Net-_C3-Pad2_ Net-_R2-Pad2_ Net-_R5-Pad2_ Net-_C1-Pad2_ Net-_Q2-Pad3_ Net-_Q2-Pad1_ Net-_C2-Pad2_ +24V Net-_C1-Pad2_ LM25085MY
R2 +24V Net-_R2-Pad2_ R
C1 +24V Net-_C1-Pad2_ CP
C2 +24V Net-_C2-Pad2_ C
C3 +24V Net-_C3-Pad2_ C
R4 +24V Net-_Q2-Pad3_ R
R3 +24V Net-_C3-Pad2_ R
D2 Net-_D2-Pad1_ Net-_C1-Pad2_ D_Schottky
Q2 Net-_Q2-Pad1_ Net-_D2-Pad1_ Net-_Q2-Pad3_ Q_PMOS_GDS
L1 Net-_D2-Pad1_ +12V L
C4 +12V Net-_C1-Pad2_ C
R5 +12V Net-_R5-Pad2_ R
R6 Net-_R5-Pad2_ Net-_C1-Pad2_ R
C5 +12V Net-_C1-Pad2_ CP
.end
