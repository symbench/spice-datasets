.title KiCad schematic
R1201 NC_01 Net-_R1201-Pad2_ Net-_R1201-Pad3_ NC_02 R_Shunt
U1201 NC_03 Net-_R1201-Pad3_ Net-_R1201-Pad2_ GND +3V3 +3V3 GND NC_04 INA240
C1201 +3V3 GND C1206
.end
