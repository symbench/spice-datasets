.title KiCad schematic
J1 CARD_1 CARD_2 CARD_3 CARD_4 CARD_5 CARD_6 CARD_7 CARD_8 CARD_9 CARD_10 CARD_11 CARD_12 CARD_13 CARD_14 CARD_15 CARD_A CARD_B CARD_C CARD_D CARD_E CARD_F CARD_H CARD_J CARD_K CARD_L CARD_M CARD_N CARD_P CARD_R CARD_S EDGE_15
J2 CARD_1 CARD_2 CARD_3 CARD_4 CARD_5 CARD_6 CARD_7 CARD_8 CARD_9 CARD_10 CARD_11 CARD_12 CARD_13 CARD_14 CARD_15 CARD_A CARD_B CARD_C CARD_D CARD_E CARD_F CARD_H CARD_J CARD_K CARD_L CARD_M CARD_N CARD_P CARD_R CARD_S EDGE_15
.end
