.title KiCad schematic
AJ2 JOY_GND JOY_GND Net-_AJ2-PadL_ NC_01 Net-_AJ2-PadR_ NC_02 AUDIO-CONNECTOR-6P-SMD-3440030P1
C8 Net-_AJ2-PadL_ JOY_GND 4700pF
R45 Net-_AJ2-PadL_ NC_03 3.3K
C9 Net-_AJ2-PadR_ JOY_GND 4700pF
R46 Net-_AJ2-PadR_ NC_04 3.3K
.end
