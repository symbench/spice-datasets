.title KiCad schematic
J2 Net-_J1-Pad4_ Net-_J1-Pad3_ Net-_J1-Pad2_ Net-_C1-Pad1_ Net-_C1-Pad2_ Net-_C4-Pad2_ Net-_J2-Pad7_ Net-_C3-Pad1_ TDA1543
J1 Net-_C1-Pad1_ Net-_J1-Pad2_ Net-_J1-Pad3_ Net-_J1-Pad4_ Net-_C1-Pad2_ Conn_01x05
C2 Net-_C1-Pad1_ Net-_C1-Pad2_ C_Small
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ C_Small
R2 Net-_C1-Pad1_ Net-_C3-Pad1_ R_Small
R3 Net-_C1-Pad1_ Net-_C4-Pad2_ R_Small
R1 Net-_C1-Pad1_ Net-_J2-Pad7_ R_Small
C3 Net-_C3-Pad1_ Net-_C3-Pad2_ C_Small
C4 Net-_C4-Pad1_ Net-_C4-Pad2_ C_Small
R5 Net-_C1-Pad1_ Net-_C4-Pad1_ R_Small
R4 Net-_C3-Pad2_ Net-_C1-Pad1_ R_Small
J3 Net-_C3-Pad2_ Net-_C1-Pad1_ Net-_C4-Pad1_ Conn_01x03
.end
