.title KiCad schematic
H1 GND MountingHole_Pad
H2 GND MountingHole_Pad
.end
