.title KiCad schematic
J1 GND GND GND GND +12V_BUS +12V_BUS +12V_BUS +5V_BUS +5V_BUS +12V_BUS Conn_02x05_Top_Bottom
J2 GND GND GND GND +12V_BUS +12V_BUS +12V_BUS +5V_BUS +5V_BUS +12V_BUS Conn_02x05_Top_Bottom
J3 GND GND GND GND +12V_BUS +12V_BUS +12V_BUS +5V_BUS +5V_BUS +12V_BUS Conn_02x05_Top_Bottom
J4 GND GND GND GND +12V_BUS +12V_BUS +12V_BUS +5V_BUS +5V_BUS +12V_BUS Conn_02x05_Top_Bottom
C9 +12V_BUS GND 100uF
C13 +12V_BUS GND 100uF
C1 +12V_BUS GND 100uF
C5 +12V_BUS GND 100uF
C2 +12V_BUS GND 100pF
C6 +12V_BUS GND 100pF
C10 +12V_BUS GND 100pF
C14 +12V_BUS GND 100pF
C11 +5V_BUS GND 100uF
C15 +5V_BUS GND 100uF
C3 +5V_BUS GND 100uF
C7 +5V_BUS GND 100uF
C4 +5V_BUS GND 100pF
C8 +5V_BUS GND 100pF
C12 +5V_BUS GND 100pF
C16 +5V_BUS GND 100pF
.end
