.title KiCad schematic
U1 Net-_RP1-Pad8_ Net-_RP1-Pad7_ Net-_RP1-Pad6_ GND SDA SCL GND +3V3 AT24C02
RP2 SCL SDA NC_01 NC_02 +3V3 +3V3 +3V3 +3V3 R_PACK4
U3 Net-_JP1-Pad2_ NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 /MUX0 /MUX1 GND /MUX3 /MUX2 Net-_R4-Pad1_ NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 +3V3 CD74HC4067SM
JP2 GND Net-_JP1-Pad2_ SolderJumper_2_Open
JP1 +3V3 Net-_JP1-Pad2_ SolderJumper_2_Bridged
RP1 +3V3 +3V3 +3V3 NC_19 NC_20 Net-_RP1-Pad6_ Net-_RP1-Pad7_ Net-_RP1-Pad8_ R_PACK4
C2 GND +3V3 C_Small
R4 Net-_R4-Pad1_ GND 10K
J1 +5V GND +3V3 NC_21 NC_22 NC_23 SDA SCL NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 /MUX3 /MUX2 /MUX0 /MUX1 GND +3V3 /MOUSE_X /MOUSE_Y /BOOT_SWITCH NC_36 Conn_01x30
J6 GND +3V3 /MOUSE_X /MOUSE_Y Conn_01x04
SW14 +3V3 /BOOT_SWITCH GND SW_SPDT
.end
