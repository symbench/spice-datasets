.title KiCad schematic
C1 +5V GND 10u
J1 /SPORT GND /VBAT /HEART_BEAT /PXX_OUT NC_01 NC_02 NC_03 Conn_JR
C2 +3V3 GND 10u
C3 +3V3 GND 100u
U3 GND +3V3 +3V3 IO36=SW_DOWN IO39=SW_RIGHT IO34=DIO0 IO35=VCC_ADC IO32=HEARTBEAT IO33=SW_LEFT IO25=SCREEN_SDA IO26=SCREEN_SCL IO27=PXX_OUT_INV IO14=SPORT IO12=SW_UP GND IO13=RST NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 IO15=DIO3 IO2=DIO2 IO0=SW_PUSH IO4=DIO1 IO16=RGBLED IO17=BUZZER IO5=SCK IO18=MISO IO19=MOSI NC_10 IO21=NSS RX0 TX0 IO22=TXEN IO23=RXEN GND GND ESP32-WROOM
J4 GND +3V3 IO26=SCREEN_SCL IO25=SCREEN_SDA Screen
U2 GND +3V3 +5V AMS1117-3.3
D5 /LED_RGB_5V NC_11 GND IO16=RGBLED WS2812B
R8 +5V /LED_RGB_5V 75
C4 /LED_RGB_5V GND 100n
U4 GND NC_12 NC_13 IO15=DIO3 IO2=DIO2 IO4=DIO1 IO34=DIO0 IO13=RST GND GND +5V IO5=SCK IO18=MISO IO19=MOSI IO21=NSS IO22=TXEN IO23=RXEN GND /ANT GND GND GND E19-XXXM30S
J3 GND TX0 RX0 Programming
AE1 /ANT GND Antenna_Dipole
Q1 /PXX_OUT GND IO27=PXX_OUT_INV BSS138
R1 +3V3 IO27=PXX_OUT_INV 1k
SW1 IO12=SW_UP IO0=SW_PUSH IO33=SW_LEFT IO39=SW_RIGHT GND IO36=SW_DOWN K1-5203UA-02
BZ1 +3V3 Net-_BZ1-Pad2_ KLJ-7525-3627
Q3 IO17=BUZZER GND Net-_BZ1-Pad2_ BSS138
R4 +3V3 IO36=SW_DOWN 10k
U1 +5V GND GND VCC MATEK_MBEC6S
R5 +3V3 IO39=SW_RIGHT 10k
D1 VCC /VBAT SS34
D2 VCC /EXT_VBAT SS34
R6 VCC IO35=VCC_ADC 10k
R7 IO35=VCC_ADC GND 1k
J2 GND /EXT_VBAT Battery
J5 GND +5V /SPORT /PXX_OUT Conn_EXT_RX
D4 IO14=SPORT GND BZT52C3V3S
R3 IO14=SPORT /SPORT 1k
R2 Net-_Q2-Pad3_ /HEART_BEAT 1k
D3 +3V3 IO14=SPORT BAT54WS
Q2 IO32=HEARTBEAT GND Net-_Q2-Pad3_ BSS138
.end
