.title KiCad schematic
U2 GND Net-_U2-Pad2_ Net-_U2-Pad2_ GND GND /LESENSE1 /LESENSE2 /LESENSE3 /LESENSE4 /LESENSE5 /LESENSE6 /LESENSE7 /USART0_TX /USART0_RX NC_01 NC_02 /USART0_CTS /USART0_RTS NC_03 GND NC_04 +3V3 NC_05 +3V3 NC_06 NC_07 NC_08 NC_09 /SWO NC_10 GND NC_11 NC_12 /SWCLK /SWDIO NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 /~nRESET GND GND GND GND GND GND GND BGM13S
R3 +3V3 Net-_R3-Pad2_ 1k
D1 GND /D- /D+ +5V SP0503BAHT
C6 +3V3 GND 4.7u
C5 +3V3 GND 0.1u
U3 NC_21 NC_22 GND /D+ /D- +3V3 +3V3 Net-_R4-Pad1_ Net-_R3-Pad2_ NC_23 NC_24 GND NC_25 NC_26 /USART0_RTS /USART0_CTS /USART0_TX /USART0_RX NC_27 NC_28 GND CP2102N-A01-GQFN20
R5 GND Net-_R4-Pad1_ 47.5k
R4 Net-_R4-Pad1_ +5V 22.1k
C1 /~nRESET GND 0.1u
U1 +5V GND +5V NC_29 +3V3 LP5907MFX-3.3
C2 +5V GND 1u
C3 +3V3 GND 1u
J2 +3V3 /SWDIO GND /SWCLK GND /SWO NC_30 NC_31 NC_32 /~nRESET Cortex SWD Connector
SW1 /~nRESET GND SW_Push
TP2 +3V3 +3.3V
TP1 +5V +5V
TP3 GND GND
C4 /LESENSE1 /LESENSE2 /LESENSE3 /LESENSE4 /LESENSE5 /LESENSE6 /LESENSE7 CapSense_01x07
J1 +5V /D- /D+ NC_33 GND GND USB_B_Micro
.end
