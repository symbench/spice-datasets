.title KiCad schematic
R1 /EXT_5V Net-_D1-Pad2_ 2kR
D1 GND Net-_D1-Pad2_ RED LED
C2 /EXT_5V GND 22uF
U1 GND +3V3 /EXT_5V AMS1117-3.3
C4 +3V3 GND 22uF
U3 GND +3V3 /EN /SENSOR_VP /SENSOR_VN /IO34 /IO35 /IO32 /IO33 /IO25 /IO26 /IO27 /IO14 /IO12 GND /IO13 /SD2 /SD3 /CMD /CLK /SD0 /SD1 /IO15 /IO2 /IO0 /IO4 /IO16 /IO17 /IO5 /IO18 /IO19 NC_01 /IO21 /RXD0 /TXD0 /IO22 /IO23 GND GND ESP32-WROOM-32
R10 +3V3 /EN 10kR
C7 /EN GND 0.1uF
C9 +3V3 GND 0.1uF
C8 +3V3 GND 22uF
C1 GND /IO0 0.1uF
SW1 GND /IO0 BOOT
C3 GND /EN 0.1uF
SW2 GND /EN EN
J2 +3V3 /EN /SENSOR_VP /SENSOR_VN /IO34 /IO35 /IO32 /IO33 /IO25 /IO26 /IO27 /IO14 /IO12 GND /IO13 /SD2 /SD3 /CMD /EXT_5V Conn_01x19
J3 GND /IO23 /IO22 /TXD0 /RXD0 /IO21 GND /IO19 /IO18 /IO5 /IO17 /IO16 /IO4 /IO0 /IO2 /IO15 /SD1 /SD0 /CLK Conn_01x19
U2 NC_02 NC_03 GND Net-_J1-Pad3_ Net-_J1-Pad2_ +3V3 +3V3 /VBUS_IC Net-_R6-Pad2_ NC_04 Net-_R9-Pad1_ NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 /RTS Net-_R7-Pad1_ Net-_R8-Pad1_ /DTR NC_17 GND CP2102N-A01-GQFN28
J1 /VBUS Net-_J1-Pad2_ Net-_J1-Pad3_ NC_18 GND GND USB_B_Micro
D2 /EXT_5V /VBUS D_Schottky
R7 Net-_R7-Pad1_ /RXD0 0R
R8 Net-_R8-Pad1_ /TXD0 0R
Q1 /RTS Net-_Q1-Pad2_ /EN S8050
Q2 /DTR Net-_Q2-Pad2_ /IO0 S8050
R2 /DTR Net-_Q1-Pad2_ 10kR
R3 /RTS Net-_Q2-Pad2_ 10kR
C5 +3V3 GND 4.7uF
C6 +3V3 GND 0.1uF
R9 Net-_R9-Pad1_ GND 10K
R6 +3V3 Net-_R6-Pad2_ 2K
R4 /VBUS /VBUS_IC 22.1K
R5 /VBUS_IC GND 47.5K
.end
