.title KiCad schematic
TP1 NC_01 TestPoint
.end
