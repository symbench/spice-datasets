.title KiCad schematic
J2 RST V0 V1 V2 V4 V3 NC_01 SDA SCL GND VDD VOUT CAP2N CAP2P CAP1P CAP1N VR NC_02 Conn_02x09_Odd_Even
R4 VDD SDA 10K
R2 VDD SCL 10K
D1 VOUT GND 8V
C2 GND VOUT 1uF
C5 CAP2P CAP2N 1uF
C8 CAP1P CAP1N 1uF
R1 VOUT GND 1M
R3 VR GND 100K
R5 VDD RST 10K
C1 GND V0 1uF
R6 V1 V2 100K
C3 GND V1 1uF
C6 GND V2 1uF
C7 V4 GND 1uF
C4 V3 GND 1uF
RV1 VR V0 NC_03 POT
R7 V3 V4 100K
Q1 Net-_Q1-Pad1_ GND BL- BC847
R8 Net-_Q1-Pad1_ BL 1K
R9 Net-_Q1-Pad1_ GND 10K
J1 VDD GND SCL SDA BL RST Conn_01x06
J3 VDD BL- Conn_01x02
C9 VDD GND 1uF
.end
