.title KiCad schematic
C1 Net-_C1-Pad1_ NC_01 1000p
L1 Output Net-_C1-Pad1_ 10u
R1 Output GND 330
P1 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 CONN_01X19
.end
