.title KiCad schematic
VR1 +24V GND Net-_FB1-Pad2_ Wurth-FDSM
F1 +24V Net-_D1-Pad1_ Fuse
D1 Net-_D1-Pad1_ NC_01 D_Schottky
D2 +24V GND D_TVS
C1 +24V GND 1u
C2 +5V GND 1u
C3 +5V GND 100n
FB1 +5V Net-_FB1-Pad2_ Ferrite_Bead
D4 Net-_D4-Pad1_ +5V RED
R1 Net-_D4-Pad1_ GND 510
D3 +5V GND D_TVS
VR2 /Wurth LED driver/LED+ /Wurth LED driver/LED+ NC_02 GND NC_03 GND /Wurth LED driver/LED- Wurth-LDHM
C4 /Wurth LED driver/LED+ /Wurth LED driver/LED- 2.2u
C5 /Wurth LED driver/LED+ GND 2.2u
C6 GND +3V3 100n
U1 NC_04 GND +3V3 NC_05 GND NC_06 NC_07 GND SN65HVD233
U2 +5V GND +5V NC_08 +3V3 ADP150AUJZ-3.3-R7
C8 +3V3 GND 100n
C7 +3V3 GND 1u
U3 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 /STM32F091/~reset NC_15 NC_16 NC_17 NC_18 GND +3V3 NC_19 NC_20 NC_21 NC_22 GND +3V3 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 GND +3V3 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 NC_43 NC_44 NC_45 NC_46 /STM32F091/swdio GND +3V3 /STM32F091/swdclk NC_47 NC_48 NC_49 NC_50 NC_51 NC_52 NC_53 NC_54 NC_55 NC_56 NC_57 NC_58 NC_59 GND +3V3 STM32F091RCTx
C17 /STM32F091/~reset GND 100n
C9 +3V3 GND 100n
C10 +3V3 GND 100n
C11 +3V3 GND 100n
C12 +3V3 GND 100n
C13 +3V3 GND 10n
C14 +3V3 GND 4.7u
C15 +3V3 GND 4.7u
C16 +3V3 GND 1u
J1 +3V3 /STM32F091/swdio GND /STM32F091/swdclk GND NC_60 NC_61 NC_62 GND /STM32F091/~reset ARM_JTAG_SWD_10
.end
