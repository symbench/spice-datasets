.title KiCad schematic
J1 VCC /BB /VCC_SENSE GND CONN_04LOCK
U1 /ISEN /COMP /FB GND GND /DR /FA /VIN LM3488QMM_NOPBDGK8-M
L1 /BB /VOUT /VIN3 GND INDUCTOR_DUAL
COUT3 5V GND 47uF
COUT1 5V GND 47uF
COUT2 5V GND 47uF
CCOMP1 /COMP GND 15nF
RFB1 /FB 5V 29.4K
CFILT1 /ISEN GND 1.5nF
RSENSE1 GND /SOURCE 0.009
CCOMP2 Net-_CCOMP2-Pad1_ GND 0.47uF
CSEP1 /VOUT /VIN3 3.3uF
CSEP2 /VOUT /VIN3 3.3uF
RFB2 GND /FB 10k
CBP1 /VIN GND 0.1uF
RFILT1 /SOURCE /ISEN 100
RFADJ1 GND /FA 76.8K
RBP1 /VIN /BB 20
RCOMP1 Net-_CCOMP2-Pad1_ /COMP 215
M1 /SOURCE /SOURCE /SOURCE /DR /VIN3 /VIN3 /VIN3 /VIN3 MOSFET_NSI4778DY
D1 5V /VOUT SL44-E3_57TDIODE_DO214AB-M
CIN1 /BB GND 3.3uF
CIN2 /BB GND 3.3uF
TP1 VCC Charger+
J2 5V GND 5V GND 5V GND 5V GND 5V GND 5V GND 5V GND NC_01 GND NC_02 NC_03 /VCC_SENSE /STAT 2X10-2MMSMD
TP2-STAT1 /STAT Charger+
.end
