.title KiCad schematic
ARDUINO1 NC_01 NC_02 NC_03 GND /E0A /E1A /E0S /E1S /E0B /E1B /LED /IN1_SENSE Net-_ARDUINO1-Pad13_ /MOSI /MISO /SCK NC_04 NC_05 Net-_ARDUINO1-Pad19_ Net-_ARDUINO1-Pad20_ Net-_ARDUINO1-Pad21_ Net-_ARDUINO1-Pad22_ /SDA /SCL NC_06 /VSENSE VCC NC_07 GND +9V ARDUINO_NANO
C2 /E1B GND 10n
C3 /E1A GND 10n
C4 /E0B GND 10n
C5 /E0A GND 10n
C6 /E0S GND 10n
C1 /E1S GND 10n
R1 VCC /SCL 3K
R2 VCC /SDA 3K
J1 GND /E0S /E0B /E0A Enc_MAIN
J2 GND /E1S /E1B /E1A Enc_INPUT
J3 GND VCC Net-_J3-Pad3_ LED
R3 Net-_J10-Pad1_ /VSENSE 510K
R4 /VSENSE GND 100K
J10 Net-_J10-Pad1_ VBAT
J14 GND +9V PWR
J11 GND /SDA /SCL Audio
J12 GND VCC /SDA /SCL LCD
C8 +9V GND 10uf
C7 +9V GND 10uf
J5 Net-_ARDUINO1-Pad22_ A3
J6 Net-_ARDUINO1-Pad21_ A2
J7 Net-_ARDUINO1-Pad20_ A1
J8 Net-_ARDUINO1-Pad19_ A0
J4 Net-_ARDUINO1-Pad13_ D10
J9 GND /SCK /MISO /MOSI SPI
J13 GND /SDA /SCL D_Pots
J15 /IN1_SENSE IN1_SENS
R5 Net-_J3-Pad3_ /LED 470
J16 GND VCC 5V
.end
