.title KiCad schematic
C86 NC_01 Net-_C86-Pad2_ C
C88 NC_02 Net-_C86-Pad2_ C
C87 Net-_C87-Pad1_ NC_03 C
C89 Net-_C87-Pad1_ NC_04 C
J32 Net-_C86-Pad2_ NC_05 Net-_J32-Pad3_ Net-_J32-Pad4_ NC_06 Net-_C87-Pad1_ InConnector
J33 NC_07 NC_08 Net-_C248-Pad1_ Net-_C249-Pad1_ NC_09 NC_10 OutConnector
C91 Net-_C249-Pad1_ NC_11 C
R239 Net-_C249-Pad1_ Net-_J32-Pad4_ R
L3 Net-_C249-Pad1_ NC_12 L
C90 Net-_C248-Pad1_ NC_13 C
R238 Net-_C248-Pad1_ Net-_J32-Pad3_ R
L2 Net-_C248-Pad1_ NC_14 L
C248 Net-_C248-Pad1_ NC_15 C
C250 Net-_C248-Pad1_ NC_16 C
C249 Net-_C249-Pad1_ NC_17 C
C251 Net-_C249-Pad1_ NC_18 C
.end
