.title KiCad schematic
U3 NC_01 /HSS_08 /HSS_07 /HSS_06 /HSS_05 /HSS_04 /HSS_03 /HSS_02 /HSS_01 /HSS_14 /HSS_13 /HSS_12 /HSS_11 /HSS_10 /HSS_09 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 IVL2-7_5
U1 /GPB7 /GPB6 /GPB5 /GPB4 /GPB3 /GPB2 /GPB1 /GPB0 +24V GND /HSS_08 /HSS_07 /HSS_06 /HSS_05 /HSS_04 /HSS_03 /HSS_02 /HSS_01 TBD62783A
U2 /GPA5 /GPA4 /GPA3 /GPA2 /GPA1 /GPA0 NC_10 NC_11 +24V GND NC_12 NC_13 /HSS_14 /HSS_13 /HSS_12 /HSS_11 /HSS_10 /HSS_09 TBD62783A
U7 /GPB0 /GPB1 /GPB2 /GPB3 /GPB4 /GPB5 /GPB6 /GPB7 +3V3 GND NC_14 NC_15 NC_16 NC_17 GND GND GND /IO_RESET NC_18 NC_19 /GPA0 /GPA1 /GPA2 /GPA3 /GPA4 /GPA5 NC_20 NC_21 MCP23017_SS
R1 +3V3 /IO_RESET 10k
.end
