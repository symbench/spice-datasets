.title KiCad schematic
U1 NC_01 NC_02 RST GND NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 LSERVO RSERVO NC_10 NC_11 TAIL NC_12 NC_13 BUZZ SENS NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 5V NC_20 GND VCC ArduinoNano
P4 GND 5V RSERVO CONN_01X03
P3 GND 5V LSERVO CONN_01X03
P1 GND Net-_P1-Pad2_ CONN_01X02
P2 GND Net-_P2-Pad2_ CONN_01X02
R2 Net-_P2-Pad2_ TAIL R
D1 Net-_D1-Pad1_ 5V LED
R1 Net-_D1-Pad1_ GND R
F1 Net-_F1-Pad1_ VCC F_Small
SW2 NC_21 Net-_P1-Pad2_ Net-_F1-Pad1_ Switch_SPDT_x2
SP1 5V Net-_D2-Pad2_ SPEAKER
SW1 RST GND SW_PUSH_SMALL_H
P5 GND 5V SENS CONN_01X03
D2 Net-_D2-Pad1_ Net-_D2-Pad2_ D
R3 5V Net-_D2-Pad1_ R
R4 Net-_Q1-Pad1_ BUZZ R
Q1 Net-_Q1-Pad1_ GND Net-_D2-Pad2_ MMBT3904
.end
