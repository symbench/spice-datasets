.title KiCad schematic
C2 +3V3 GND 100nF
J1 +3V3 /SDA /SCL /GP4 GND I2C
C1 +3V3 GND 100nF
J4 GND +3V3 /SDA /SCL GND QWIIC1
J6 GND +3V3 /SDA /SCL GND QWIIC2
J3 /MOSI /MISO Net-_J3-Pad3_ /CS +3V3 GND Net-_J3-Pad7_ /PCM_DIN /PCM_DOUT /PCM_FS GND +5V SPI_I2S
J5 +3V3 +5V /SDA +5V /SCL GND /GP4 Net-_J2-Pad8_ GND Net-_J2-Pad10_ Net-_J2-Pad11_ Net-_J2-Pad12_ Net-_J2-Pad13_ GND Net-_J2-Pad15_ Net-_J2-Pad16_ +3V3 /PCM_CLK /MOSI GND /MISO Net-_J2-Pad22_ /SCK /CS0 GND /CS1 Net-_J2-Pad27_ Net-_J2-Pad28_ Net-_J2-Pad29_ GND Net-_J2-Pad31_ Net-_J2-Pad32_ Net-_J2-Pad33_ GND /PCM_FS Net-_J2-Pad36_ Net-_J2-Pad37_ /PCM_DIN GND /PCM_DOUT RPI_IN
J2 +3V3 +5V /SDA +5V /SCL GND /GP4 Net-_J2-Pad8_ GND Net-_J2-Pad10_ Net-_J2-Pad11_ Net-_J2-Pad12_ Net-_J2-Pad13_ GND Net-_J2-Pad15_ Net-_J2-Pad16_ +3V3 /PCM_CLK /MOSI GND /MISO Net-_J2-Pad22_ /SCK /CS0 GND /CS1 Net-_J2-Pad27_ Net-_J2-Pad28_ Net-_J2-Pad29_ GND Net-_J2-Pad31_ Net-_J2-Pad32_ Net-_J2-Pad33_ GND /PCM_FS Net-_J2-Pad36_ Net-_J2-Pad37_ /PCM_DIN GND /PCM_DOUT RPI_IN
JP1 /CS0 /CS /CS1 SPI CS
C4 +5V GND 100nF
C3 +3V3 GND 100nF
R1 /SCK Net-_J3-Pad3_ 47R
R2 /PCM_CLK Net-_J3-Pad7_ 47R
.end
