.title KiCad schematic
U1 Net-_R7-Pad1_ Net-_C5-Pad1_ Net-_C5-Pad1_ NC_01 ~SHORT Net-_C5-Pad1_ NC_02 NC_03 EN/UVLO IVINP IVINN Vin INTVcc1 TG1 BST1 SW1 SNSN1 BG1 BG2 SNSN1 SW2 BST2 NC_04 TG2 ISP ISN SNSP1 SNSN1 NC_05 SNSN1 NC_06 INTVcc1 NC_07 SNSN1 Net-_R11-Pad2_ Net-_R9-Pad2_ FB OVLO LT3790
Q1 SW1 SW1 SW1 TG1 Vin Vin Vin Vin BSC123N10LSGATMA1
R7 Net-_R7-Pad1_ Net-_C5-Pad1_ R
C5 Net-_C5-Pad1_ SNSN1 33n
R8 INTVcc1 ~SHORT 200k
C6 SNSN1 Net-_C5-Pad1_ 100n
R5 IVINP OVLO 150k
R6 OVLO SNSN1 10k
R3 IVINP EN/UVLO 10k
R4 EN/UVLO SNSN1 20k
C2 EN/UVLO SNSN1 220p
R9 Net-_C8-Pad2_ Net-_R9-Pad2_ 3,3k
C8 SNSN1 Net-_C8-Pad2_ 33n
R1 Vin IVINP 3m
C1 IVINN IVINP 470n
C3 Vin SNSN1 4.7u
C4 Vin SNSN1 4.7u
C7 Vin SNSN1 1u
R2 Vin IVINN 51
D2 BST1 INTVcc1 D_Schottky
C10 BST1 SW1 100n
Q2 SNSP1 SNSP1 SNSP1 BG1 SW1 SW1 SW1 SW1 BSC123N10LSGATMA1
R10 SNSP1 SNSN1 4m
Q3 SW2 SW2 SW2 TG2 ISP ISP ISP ISP BSC123N10LSGATMA1
C11 BST2 SW2 100n
Q4 SNSP1 SNSP1 SNSP1 BG2 SW2 SW2 SW2 SW2 BSC123N10LSGATMA1
L1 SW2 SW1 10u
R12 PWR_OUT ISP 4m
C12 ISP SNSN1 4.7u
R13 PWR_OUT ISN 51
C13 ISN ISP 0.47u
C9 INTVcc1 SNSN1 100n
C14 PWR_OUT SNSN1 220u
R14 FB PWR_OUT 58k
R15 SNSN1 FB 1.2k
R11 SNSN1 Net-_R11-Pad2_ 147k
D1 BST2 INTVcc1 D_Schottky
.end
