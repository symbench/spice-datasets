.title KiCad schematic
J1 /RGB4 /RGB3 /RGB2 /RGB1 /RGB0 Conn_01x05
J2 /ROW0 /ROW1 /ROW2 /ROW3 /ROW4 Conn_01x05
J3 /MUX3 /MUX2 /MUX0 /MUX1 Conn_01x04
J4 GND /USB_D- /USB_D+ +5V Conn_01x04
J5 GND GND GND GND GND Conn_01x05
J6 +3V3 +3V3 +3V3 +3V3 +3V3 Conn_01x05
J7 /SDA /SCL Conn_01x02
J8 /LED0 /LED1 /LED2 Conn_01x03
J11 +5V GND +3V3 /LED0 /LED1 /LED2 /SDA /SCL /USB_D- /USB_D+ /RGB4 /RGB3 /RGB2 /RGB1 /RGB0 /ROW0 /ROW1 /ROW2 /ROW3 /ROW4 /MUX3 /MUX2 /MUX0 /MUX1 GND +3V3 /MOUSE_X /MOUSE_Y /BOOT_SWITCH NC_01 Conn_01x30
J12 +5V GND +3V3 /LED0 /LED1 /LED2 /SDA /SCL /USB_D- /USB_D+ /RGB4 /RGB3 /RGB2 /RGB1 /RGB0 /ROW0 /ROW1 /ROW2 /ROW3 /ROW4 /MUX3 /MUX2 /MUX0 /MUX1 GND +3V3 /MOUSE_X /MOUSE_Y /BOOT_SWITCH NC_02 Conn_01x30
J9 /MOUSE_X /MOUSE_Y GND Conn_01x03
J10 /BOOT_SWITCH GND Conn_01x02
.end
