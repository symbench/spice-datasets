.title KiCad schematic
LOGO1 BUTTERFLY_LOGO
R9 GND SW_FUNCTION 47K
R10 GND SW_SELECT 47K
R17 GND SW_RESET 47K
R44 Net-_LED4-PadA_ /LED4 390
R43 Net-_LED3-PadA_ /LED3 390
R27 Net-_LED2-PadA_ /LED2 390
R26 Net-_LED1-PadA_ /LED1 390
LED4 Net-_LED4-PadA_ GND LEDCHIPLED_0603
LED3 Net-_LED3-PadA_ GND LEDCHIPLED_0603
LED2 Net-_LED2-PadA_ GND LEDCHIPLED_0603
LED1 Net-_LED1-PadA_ GND LEDCHIPLED_0603
S3 SW_FUNCTION SW_FUNCTION 3V3_PWR6 3V3_PWR6 EVQQ2
S1 SW_SELECT SW_SELECT 3V3_PWR6 3V3_PWR6 EVQQ2
S4 SW_RESET SW_RESET 3V3_PWR6 3V3_PWR6 EVQQ2
H1 3V3_PWR6 5V0 5V 5V NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 SW_SELECT NC_27 SW_RESET NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 /PS2CLK2 NC_36 /PS2DAT2 NC_37 NC_38 NC_39 NC_40 NC_41 /LED1 NC_42 /LED2 NC_43 /LED3 NC_44 /LED4 GND GND GND GND GND NC_45 NC_46 NC_47 NC_48 Arduino Mega Header
PWR_2 GND NC_49 3V3_PWR6 5V0 POWER_ONLYNOTEXT
PWR_1 GND NC_50 3V3_PWR6 NC_51 POWER_ONLYNOTEXT
R47 /PS2DAT2 Net-_PS2_B1-Pad1_ 390
R48 /PS2CLK2 Net-_PS2_B1-Pad5_ 390
PS2_B1 Net-_PS2_B1-Pad1_ NC_52 GND 5V0 Net-_PS2_B1-Pad5_ NC_53 MINI-DIN6PTH
.end
