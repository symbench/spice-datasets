.title KiCad schematic
IC1 Net-_IC1-Pad1_ NC_01 NC_02 Net-_IC1-Pad4_ Net-_IC1-Pad5_ Net-_IC1-Pad6_ Net-_IC1-Pad7_ /BUFFEN Net-_IC1-Pad9_ GND Net-_IC1-Pad11_ Net-_IC1-Pad12_ NC_03 NC_04 NC_05 /RST /MOSI /MISO /SCK VCC ATTINY2313-S
U2 /BUFFEN /SCK Net-_R1-Pad2_ /BUFFEN /RST /RST' GND Net-_R2-Pad2_ /MOSI /BUFFEN /MISO /MISO' /BUFFEN VCC 74LS125
X1 Net-_IC1-Pad4_ Net-_IC1-Pad5_ GND CRYSTAL_SMD
P2 VCC Net-_D4-Pad1_ Net-_D3-Pad1_ GND GND GND USB_OTG
C1 VCC GND 100U
R3 Net-_D3-Pad1_ Net-_IC1-Pad6_ 47
R6 Net-_D4-Pad1_ Net-_IC1-Pad7_ 47
D2 GND Net-_D2-Pad2_ LED
D1 GND Net-_D1-Pad2_ LED
R7 Net-_D2-Pad2_ Net-_IC1-Pad12_ 1K
R4 Net-_D1-Pad2_ Net-_IC1-Pad9_ 1K
P1 /MISO' VCC /SCK' /MOSI' /RST' GND CONN_02X03
R2 /MOSI' Net-_R2-Pad2_ 1.5K
R1 /SCK' Net-_R1-Pad2_ 1.5K
C2 VCC GND 0.1U
D3 Net-_D3-Pad1_ GND D
D4 Net-_D4-Pad1_ GND D
R5 Net-_D4-Pad1_ Net-_IC1-Pad11_ 1.5K
P3 /MISO VCC /SCK /MOSI /RST GND CONN_02X03
R8 Net-_IC1-Pad1_ VCC 10K
.end
