.title KiCad schematic
U1 VCC GND VCC Net-_C1-Pad1_ +3V3 MIC5219-3.3
J1 GND VCC PA10=RX PA9=TX Conn_01x04_Female
J2 GND SWCLK SWDIO +3V3 Conn_01x04_Female
C1 Net-_C1-Pad1_ GND 470p
C2 +3V3 GND 2.2u
C3 +3V3 GND 100n
C4 +3V3 GND 100n
C5 +3V3 GND 100n
C6 +3V3 GND 100n
Y1 Net-_U2-Pad5_ GND Net-_U2-Pad6_ 8Mhz
U2 +3V3 NC_01 NC_02 NC_03 Net-_U2-Pad5_ Net-_U2-Pad6_ +3V3 GND +3V3 NC_04 NC_05 NC_06 NC_07 PA4=NSS PA5=SCK PA6=MISO PA7=MOSI PB0=NRESET PB1=BUSY NC_08 PB10=DIO1 PB11=LED GND +3V3 NC_09 NC_10 NC_11 NC_12 NC_13 PA9=TX PA10=RX Net-_SW1-Pad1_ NC_14 SWDIO GND +3V3 SWCLK NC_15 NC_16 PB4=RX_EN PB5=TX_EN PB6=DIO2 NC_17 GND NC_18 NC_19 GND +3V3 STM32F103C8Tx
D1 GND Net-_D1-Pad2_ LED
R1 PB11=LED Net-_D1-Pad2_ R
SW1 Net-_SW1-Pad1_ GND SW_Push
U3 GND GND GND GND GND PB4=RX_EN PB5=TX_EN PB6=DIO2 +3V3 GND GND GND PB10=DIO1 PB1=BUSY PB0=NRESET PA6=MISO PA7=MOSI PA5=SCK PA4=NSS GND NC_20 GND E22-X00M22S
.end
