.title KiCad schematic
J4 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 GND NC_09 NC_10 GND NC_11 NC_12 NC_13 NC_14 691327310016
J5 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 691327310016
U1 5V GND NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 NC_43 NC_44 NC_45 NC_46 NC_47 NC_48 NC_49 NC_50 NC_51 NC_52 NC_53 GND NC_54 NC_55 NC_56 NC_57 NC_58 NC_59 NC_60 NC_61 GND NC_62 5V 5V NC_63 GND GND NC_64 GND Net-_U1-Pad44_ Net-_U1-Pad44_ GND GND 5V NC_65 NC_66 NC_67 GND NC_68 GND GND GND NC_69 GND NC_70 GND NC_71 NC_72 GND GND ADS8586S
U6 NC_73 NC_74 NC_75 NC_76 NC_77 NC_78 NC_79 NC_80 THS4032ID
U8 NC_81 NC_82 5V NC_83 NC_84 GND NC_85 NC_86 THS4551IDGKT
U7 NC_87 NC_88 5V NC_89 NC_90 GND NC_91 NC_92 THS4551IDGKT
J16 NC_93 GND NC_94 NC_95 NC_96 NC_97 GND MDD01
.end
