.title KiCad schematic
J1 Net-_C3-Pad1_ /USBD- /USBD+ GND GND USB_B
F1 +5V Net-_C3-Pad1_ F_500mA_16V
C3 Net-_C3-Pad1_ GND C_100nF
U2 +5V GND +5V NC_01 +3V3 MIC5205-3.3YM5
C6 +3V3 GND C_10uF
C7 +3V3 GND C_0.1uF
C1 +5V GND C_0.1uF
C4 +5V GND C_10uF
U1 NC_02 NC_03 +5V Net-_R3-Pad2_ NC_04 GND NC_05 NC_06 NC_07 Net-_D4-Pad1_ /USBD+ /USBD- /3V3_FTDI /3V3_FTDI /3V3_FTDI GND Net-_D2-Pad1_ NC_08 NC_09 Net-_R2-Pad2_ FT231XS
C2 /3V3_FTDI GND C_0.1uF
R2 /Rx Net-_R2-Pad2_ R_1K
R3 /Tx Net-_R3-Pad2_ R_1K
U3 NC_10 NC_11 GND +5V GND +5V /XTAL1 /XTAL2 NC_12 NC_13 NC_14 /IO8 NC_15 NC_16 /MOSI /MISO /SCK +5V NC_17 /AREF GND NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 /RST /Rx /Tx NC_25 ATmega328P-AU
J3 /MISO +5V /SCK /MOSI /RST GND CONN_02X03
D2 Net-_D2-Pad1_ Net-_D2-Pad2_ LED
D4 Net-_D4-Pad1_ Net-_D4-Pad2_ LED
R7 +5V Net-_D4-Pad2_ R_1K
R6 +5V Net-_D2-Pad2_ R_1K
D1 Net-_D1-Pad1_ +5V 5V_LED
R1 Net-_D1-Pad1_ GND R_1K
D3 Net-_D3-Pad1_ +3V3 LED
R4 Net-_D3-Pad1_ GND R_1K
R5 Net-_D5-Pad1_ GND R_1K
D7 Net-_D7-Pad1_ /SCK LED
R8 Net-_D7-Pad1_ GND R_1K
D8 Net-_D8-Pad1_ /IO8 LED
R9 Net-_D8-Pad1_ GND R_1K
D6 /Vin Net-_D6-Pad2_ CDBA140-G
C8 /Vin GND C_47uF
D5 Net-_D5-Pad1_ /Vin LED
U4 GND +5V /Vin LM1117-5.0
J2 Net-_D6-Pad2_ GND Barrel_Jack
C10 +5V GND C_0.1uF
C9 +5V GND C_10uF
Y1 /XTAL1 GND /XTAL2 GND Crystal_SMD
C11 /XTAL1 GND C_30pF
C12 /XTAL2 GND C_30pF
C5 /AREF GND C_0.1uF
.end
