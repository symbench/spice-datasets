.title KiCad schematic
K2 Net-_K2-Pad1_ Net-_K2-Pad1_ Net-_K2-Pad3_ Net-_K2-Pad3_ Net-_K2-Pad5_ Net-_K2-Pad5_ NC_01 NC_02 NC_03 NC_04 NC_05 Maxon-200142
K1 Net-_K1-Pad1_ Net-_K1-Pad1_ Net-_K1-Pad3_ Net-_K1-Pad3_ Net-_K1-Pad5_ Net-_K1-Pad5_ NC_06 NC_07 NC_08 NC_09 NC_10 Maxon-200142
.end
