.title KiCad schematic
U1 NC_01 NC_02 Net-_U1-Pad3_ NC_03 NC_04 NC_05 Net-_U1-Pad3_ NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 AS5304
U2 NC_19 NC_20 Net-_U2-Pad3_ NC_21 NC_22 NC_23 Net-_U2-Pad3_ NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 AS5304
.end
