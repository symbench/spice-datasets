.title KiCad schematic
RV1 GND Net-_RV1-Pad2_ Net-_J1-PadT_ A100K
R2 CVIN Net-_J3-PadT_ 100K
RV3 -12V Net-_R3-Pad2_ +12V B50K
R3 CVIN Net-_R3-Pad2_ 100K
RV2 GND VERT Net-_J2-PadT_ A100K
R1 V2 Net-_J2-PadT_ 47K
J2 GND Net-_J2-PadT_ NC_01 CV1
J3 GND Net-_J3-PadT_ NC_02 CV2
J1 GND Net-_J1-PadT_ NC_03 IN
J5 S2 NC_04 V2 OUT VERT IN Conn_01x06
J6 GND CVIN +12V QR -12V QW Conn_01x06
J4 GND Net-_J4-PadT_ NC_05 OUT
R7 Net-_J4-PadT_ OUT 47K
RV4 GND QW QR A100K
SW1 Net-_R5-Pad2_ GND S2 S2 Net-_RV1-Pad2_ Net-_R5-Pad2_ SW_Push_DPDT
R5 IN Net-_R5-Pad2_ 68K
.end
