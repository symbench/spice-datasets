.title KiCad schematic
J1 +3V3 +3V3 GND +5V GND +5V NC_01 PWR_OK_RAW +5VSB +12V +12V +3V3 +3V3 -12V GND PS_ON GND GND GND -5V +5V +5V +5V GND ATX_24PIN
J2 GND GND GND GND +12V +12V +12V +12V ATX_EPS12V
J5 +12V +12V +12V GND GND GND ATX_PCIE_6PIN
J3 GND GND GND GND +12V +12V +12V +12V ATX_EPS12V
J6 +12V +12V +12V GND GND GND ATX_PCIE_6PIN
J7 +12V +12V +12V GND GND GND ATX_PCIE_6PIN
D1 NC_02 NC_03 LED_SB
R1 GND NC_04 470
D3 NC_05 NC_06 LED_OK
R3 GND NC_07 470
D2 NC_08 NC_09 LED_SW
R2 PS_ON NC_10 470
J4 +12V +12V +12V GND GND GND ATX_PCIE_6PIN
P3 NC_11 GND NC_12 GND NC_13 GND NC_14 GND NC_15 GND PWR_OK_BUF GND PS_ON GND NC_16 GND CONN_MISC
P4 GND +12V GND +12V GND +12V CONN_12V_1
P5 +12V GND +12V GND +12V GND CONN_12V_2
P6 GND +3V3 GND +3V3 CONN_3V3
P7 +5V GND +5V GND CONN_5V
JP4 +12V +12V JUMPER
U1 GND PWR_OK_RAW GND PWR_OK_BUF +5VSB LOGIC_BUFFER_3ST
P1 PWR_OK_RAW CONN_01X01
P2 PWR_OK_BUF CONN_01X01
.end
