.title KiCad schematic
U1 VCC GND VCC NC_01 +3V3 MIC5219-3.3
J1 GND VCC PA10=RX PA9=TX DATA
J2 GND SWCLK SWDIO +3V3 Programming
C2 +3V3 GND 1u
C3 +3V3 GND 100n
C4 +3V3 GND 100n
C5 +3V3 GND 100n
C6 +3V3 GND 100n
Y1 Net-_U2-Pad5_ GND Net-_U2-Pad6_ 8Mhz
U2 +3V3 NC_02 NC_03 NC_04 Net-_U2-Pad5_ Net-_U2-Pad6_ +3V3 GND +3V3 NC_05 NC_06 NC_07 NC_08 PA4=NSS PA5=SCK PA6=MISO PA7=MOSI PB0=RESET PB1=DIO3 NC_09 PB10=DIO5 PB11=LED GND +3V3 NC_10 NC_11 NC_12 NC_13 NC_14 PA9=TX PA10=RX Net-_SW1-Pad1_ NC_15 SWDIO GND +3V3 SWCLK NC_16 NC_17 PB4=DIO2 PB5=DIO1 PB6=DIO0 PB7=DIO4 GND PB8 PB9 GND +3V3 STM32F103C8Tx
D1 GND Net-_D1-Pad2_ LED
R1 PB11=LED Net-_D1-Pad2_ R
SW1 Net-_SW1-Pad1_ GND SW_Push
U3 GND PA6=MISO PA7=MOSI PA5=SCK PA4=NSS PB0=RESET PB10=DIO5 GND /ANT GND PB1=DIO3 PB7=DIO4 +3V3 PB6=DIO0 PB5=DIO1 PB4=DIO2 RFM95W-868S2
AE1 /ANT GND Antenna_Dipole
J3 GND PB8 PB9 +3V3 Expansion
.end
