.title KiCad schematic
U3 NC_01 Net-_U3-Pad2_ NC_02 Net-_U3-Pad2_ NC_03 NC_04 SY8105
.end
