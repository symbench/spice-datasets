.title KiCad schematic
C1 +3V3 GND 10u
C3 +3V3 GND 10n
C4 +3V3 GND 10n
C6 +3V3 GND 10n
C5 GND /NRF_XC1 22p
C7 GND /NRF_XC2 22p
R2 /NRF_XC1 /NRF_XC2 1M
C2 GND Net-_C2-Pad2_ 22p
U1 NRF_CE NC_01 NC_02 NC_03 NC_04 NC_05 +3V3 GND /NRF_XC2 /NRF_XC1 /NRF_VDD_PA /NRF_ANT1 /NRF_ANT2 GND +3V3 Net-_R1-Pad1_ GND +3V3 Net-_C2-Pad2_ GND nRF24L01P
R1 Net-_R1-Pad1_ GND 22k
C9 +3V3 GND 10n
C8 +3V3 GND 220p
C10 +3V3 GND 2u2
C11 GND /RFX_ANT 22p
J1 GND GND GND GND Net-_F1-Pad5_ 5-1814400-1
C12 /NRF_VDD_PA GND 2n2
C14 /NRF_VDD_PA GND 4p7
C15 /RFX_TXRX GND 22p
C13 Net-_C13-Pad1_ /RFX_TXRX 22p
L3 /NRF_ANT2 /NRF_VDD_PA 2n7
L2 /NRF_ANT1 Net-_C13-Pad1_ 3n9
L1 /NRF_ANT1 /NRF_ANT2 8n2
F1 GND /RFX_ANT GND GND Net-_F1-Pad5_ GND 2450LP14B100
Y1 /NRF_XC1 GND GND /NRF_XC2 16MHz
IC1 GND GND GND /RFX_TXRX /NRF_VDD_PA NRF_CE GND GND GND /RFX_ANT GND GND NC_06 +3V3 GND +3V3 GND RFX2401C
.end
