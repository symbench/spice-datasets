.title KiCad schematic
U1 NC_01 /RGB4 /RGB2 /RGB0 /LED0 /LED1 /LED2 /ROW0 /ROW1 /ROW2 /ROW3 /ROW4 /MOUSE_X /MOUSE_Y NC_02 NC_03 NC_04 +3V3 GND GND NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 /USB_D- /USB_D+ NC_12 /BOOT_SWITCH /MUX1 /MUX0 /SCL /SDA /MUX2 /MUX3 +5V GND +3V3 NC_13 NC_14 BluePill_STM32F103C
J1 +3V3 GND /MUX1 /MUX0 /MUX2 /MUX3 /ROW4 /ROW3 /ROW2 /ROW1 /ROW0 /RGB0 NC_15 /RGB2 NC_16 /RGB4 /USB_D+ /USB_D- /SCL /SDA /LED2 /LED1 /LED0 +3V3 GND +5V /MOUSE_X /MOUSE_Y /BOOT_SWITCH NC_17 Conn_01x30
.end
