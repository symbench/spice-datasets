.title KiCad schematic
U1 GND Net-_C2-Pad2_ Net-_R3-Pad2_ 5V Net-_C1-Pad2_ Net-_C2-Pad2_ Net-_R1-Pad1_ VCC LM555N
C1 GND Net-_C1-Pad2_ 10n
R2 Net-_R1-Pad1_ Net-_C2-Pad2_ 12k
R1 Net-_R1-Pad1_ 5V 2.2k
1N400X1 Net-_1N400X1-Pad1_ VCC D
C3 Net-_1N400X1-Pad1_ GND 220u
C4 12V GND 47u
C5 5V GND 47u
R5 Net-_D1-Pad2_ 5V 270
D1 GND Net-_D1-Pad2_ LED
2N1 Net-_2N1-Pad1_ Net-_2N1-Pad2_ GND Q_NPN_BCE
R4 Net-_1N400X1-Pad1_ Net-_2N1-Pad2_ 1.8k
2N2222_1 Net-_2N1-Pad2_ Net-_1N400X1-Pad1_ Net-_2N2-Pad3_ Q_NPN_BCE
2N2 Net-_2N1-Pad2_ GND Net-_2N2-Pad3_ Q_PNP_BCE
C7 Net-_2N2-Pad3_ Net-_1N400X2-Pad2_ 47u
1N400X2 GND Net-_1N400X2-Pad2_ D
1N400X3 Net-_1N400X2-Pad2_ Net-_1N400X3-Pad2_ D
C8 GND Net-_1N400X3-Pad2_ 47u
C9 GND -12V 47u
R3 Net-_2N1-Pad1_ Net-_R3-Pad2_ 3.3k
C2 GND Net-_C2-Pad2_ 47n
U5 GND Net-_1N400X3-Pad2_ -12V LM2990T-12
U6 GND -12V -5V LM2990T-5
C10 GND -5V 47u
U2 GND Net-_1N400X1-Pad1_ 12V LM2940CT-12
U3 GND 12V 5V LM2940CT-5
U4 GND 12V 3.3V LM1117T-3.3
C6 3.3V GND 47u
.end
