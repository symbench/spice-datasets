.title KiCad schematic
J1 Net-_J1-Pad1_ Net-_J1-Pad2_ Net-_J1-Pad3_ C
J2 Net-_J1-Pad1_ Net-_J1-Pad2_ Net-_J1-Pad3_ C
J3 Net-_J1-Pad1_ Net-_J1-Pad2_ Net-_J1-Pad3_ C
.end
