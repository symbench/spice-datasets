.title KiCad schematic
U1 TXD RXD VBAT +3V3 GND PPS GND GND GND GND GND GND GND SKM61
P1 PPS GND +3V3 VBAT RXD TXD CONN_01X06
.end
