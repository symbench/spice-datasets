.title KiCad schematic
IC1 /SCHW_1/MOSI/SDA /SCHW_1/MISO /SCHW_1/SCK NC_01 VCC GND NC_02 NC_03 NC_04 /SCHW_1/RESET NC_05 /SCHW_1/RIGHT /SCHW_1/ENC_A_RAW /SCHW_1/ENC_B_RAW VCC GND /SCHW_1/DOWN /SCHW_1/OK /SCHW_1/UP /SCHW_1/LEFT TINY26S
R1 /SCHW_1/RESET VCC 10k
R2 /SCHW_1/ENC_B_RAW /SCHW_1/ENC_B 10K
R3 /SCHW_1/ENC_A_RAW /SCHW_1/ENC_A 10K
C1 GND VCC 100n
C2 /SCHW_1/ENC_A GND 100n
C3 /SCHW_1/ENC_B GND 100n
BUTTONS1 /SCHW_1/ENC_A /SCHW_1/ENC_B GND GND /SCHW_1/OK /SCHW_1/DOWN /SCHW_1/RIGHT /SCHW_1/UP /SCHW_1/LEFT ENCODER_ARROWS
POWER1 VCC NC_06 PINHD-1X2
OLED1 Net-_J2-Pad2_ Net-_J1-Pad2_ /SCHW_1/SCK /SCHW_1/MOSI/SDA PINHD-1X4
PROG1 /SCHW_1/MOSI/SDA /SCHW_1/MISO /SCHW_1/SCK /SCHW_1/RESET VCC GND PINHD-1X6
J1 GND Net-_J1-Pad2_ VCC SJ2W
J2 GND Net-_J2-Pad2_ VCC SJ2W
T1 NC_07 GND NC_08 AP2306GN_MOSFETSOT23
.end
