.title KiCad schematic
U1 GND /SCL /SDA NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 /LCD_CS /SCK /MISO /MOSI NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 /LCD_BL NC_17 NC_18 /LCD_DC /LCD_RST /T_CS /T_IRQ NC_19 NC_20 +3V3 GND blackpill
J3 +3V3 GND /SCL /SDA NC_21 NC_22 Conn_01x06
J2 GND GND Conn_01x02
J1 /T_IRQ /MISO /MOSI /T_CS /SCK /MISO /LCD_BL /SCK /MOSI /LCD_DC /LCD_RST /LCD_CS GND +3V3 Conn_01x14
J4 GND +3V3 /SCK /MOSI /LCD_RST /LCD_DC /LCD_BL Conn_01x07
.end
