.title KiCad schematic
BT1 Net-_BT1-Pad1_ Net-_BT1-Pad2_ Battery_Cell
J1 Net-_BT1-Pad1_ Net-_BT1-Pad1_ Net-_BT1-Pad1_ Conn_01x03_Female
J2 Net-_BT1-Pad2_ Net-_BT1-Pad2_ Net-_BT1-Pad2_ Conn_01x03_Female
.end
