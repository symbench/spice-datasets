.title KiCad schematic
U12 +3V3 XBEE_DEBUG_EN NC_01 NC_02 GND CC_UART0_TX CC_UART0_RX XBEE_DEBUG_RX XBEE_DEBUG_TX Net-_R28-Pad2_ FSUSB42MUX
R28 GND Net-_R28-Pad2_ 10k
C48 +3V3 GND 4.7uF
C50 +3V3 GND 0.1uF
R26 GND XBEE_DEBUG_EN 10k
U11 +3V3 GPS_DEBUG_EN NC_03 NC_04 GND NC_05 NC_06 GPS_DEBUG_RX GPS_DEBUG_TX Net-_R27-Pad2_ FSUSB42MUX
R27 GND Net-_R27-Pad2_ 10k
C47 +3V3 GND 4.7uF
C49 +3V3 GND 0.1uF
R25 GND GPS_DEBUG_EN 10k
J5 NC_07 GND Conn_01x02
J1 VBUS VBUS VBUS VBUS GPS_DEBUG_EN GPS_DEBUG_RX GPS_DEBUG_TX NC_08 XBEE_DEBUG_TX XBEE_DEBUG_RX XBEE_DEBUG_EN NC_09 NC_10 NC_11 NC_12 NC_13 CC_UART0_TX CC_UART0_RX NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 +3V3 +3V3 GND GND GND GND Conn_02x18_Odd_Even
.end
