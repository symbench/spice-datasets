.title KiCad schematic
U2 GND ~BUSACK Net-_R5-Pad1_ ~BUSRQ Net-_R6-Pad1_ ~IORQ Net-_R7-Pad1_ ~MREQ Net-_R8-Pad1_ GND ~M1 Net-_R4-Pad1_ ~HALT Net-_R3-Pad1_ ~RD Net-_R2-Pad1_ ~WR Net-_R1-Pad1_ GND VCC 74HC240
R8 Net-_R8-Pad1_ Net-_M1-Pad2_ 330
R7 Net-_R7-Pad1_ Net-_HALT1-Pad2_ 330
R6 Net-_R6-Pad1_ Net-_R6-Pad2_ 330
R5 Net-_R5-Pad1_ Net-_R5-Pad2_ 330
R4 Net-_R4-Pad1_ Net-_MREQ1-Pad2_ 330
R3 Net-_R3-Pad1_ Net-_IORQ1-Pad2_ 330
R2 Net-_R2-Pad1_ Net-_BUSRQ1-Pad2_ 330
R1 Net-_R1-Pad1_ Net-_BUSACK1-Pad2_ 330
M1 GND Net-_M1-Pad2_ LED_ALT
HALT1 GND Net-_HALT1-Pad2_ LED_ALT
RD1 GND Net-_R6-Pad2_ LED_ALT
WR1 GND Net-_R5-Pad2_ LED_ALT
MREQ1 GND Net-_MREQ1-Pad2_ LED_ALT
IORQ1 GND Net-_IORQ1-Pad2_ LED_ALT
BUSRQ1 GND Net-_BUSRQ1-Pad2_ LED_ALT
BUSACK1 GND Net-_BUSACK1-Pad2_ LED_ALT
J1 ~M1 ~HALT ~RD ~WR ~MREQ ~IORQ ~BUSRQ ~BUSACK GND VCC Conn_01x10
C1 VCC GND 100 nF
.end
