.title KiCad schematic
U4 NC_01 Net-_U4-Pad2_ NC_02 Net-_U4-Pad2_ Dual_battery
.end
