.title KiCad schematic
J1 VCC DIN CLK LATCH GND RST DOUT OE 595
J2 VCC DIN CLK LATCH GND RST IN
J3 VCC DOUT CLK LATCH GND RST OUT
J4 OE OE
.end
