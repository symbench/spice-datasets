.title KiCad schematic
U1 Net-_C2-Pad1_ Net-_C3-Pad1_ GND +5V Net-_J3-Pad5_ Net-_J3-Pad3_ Net-_J3-Pad4_ RX Net-_RN3-Pad3_ Net-_RN3-Pad2_ Net-_RN3-Pad1_ Net-_J3-Pad2_ CTS NC_01 SCK MOSI MISO Net-_J4-Pad4_ Net-_J4-Pad6_ Net-_J4-Pad8_ Net-_J4-Pad10_ Net-_J4-Pad9_ Net-_J4-Pad7_ RST Net-_J4-Pad5_ Net-_J4-Pad3_ Net-_C4-Pad1_ GND Net-_RN1-Pad3_ Net-_RN1-Pad2_ +5V +5V ATMEGA8U2-AU
RN2 GND NC_02 Net-_D1-Pad1_ +5V RST GND NC_03 CTS R_Pack04
RN3 Net-_RN3-Pad1_ Net-_RN3-Pad2_ Net-_RN3-Pad3_ Net-_RN3-Pad3_ TX TX Net-_D2-Pad1_ Net-_D3-Pad1_ R_Pack04
RN1 NC_04 Net-_RN1-Pad2_ Net-_RN1-Pad3_ NC_05 NC_06 Net-_J1-Pad3_ Net-_J1-Pad2_ NC_07 22R
J1 Net-_F1-Pad2_ Net-_J1-Pad2_ Net-_J1-Pad3_ NC_08 GND GND USB_OTG
F1 +5V Net-_F1-Pad2_ Fuse
CON1 MISO +5V SCK MOSI RST GND AVR-ISP-6
Y1 Net-_C2-Pad1_ Net-_C3-Pad1_ Crystal
C2 Net-_C2-Pad1_ GND 22pF
C3 Net-_C3-Pad1_ GND 22pF
C4 Net-_C4-Pad1_ GND 1uF
D1 Net-_D1-Pad1_ +5V P
D2 Net-_D2-Pad1_ +5V R
D3 Net-_D3-Pad1_ +5V T
J2 CTS RX TX +5V GND GND Conn_01x06
C1 +5V GND 100n
C5 +5V GND 100n
J4 +5V GND Net-_J4-Pad3_ Net-_J4-Pad4_ Net-_J4-Pad5_ Net-_J4-Pad6_ Net-_J4-Pad7_ Net-_J4-Pad8_ Net-_J4-Pad9_ Net-_J4-Pad10_ EXP1
J3 +5V Net-_J3-Pad2_ Net-_J3-Pad3_ Net-_J3-Pad4_ Net-_J3-Pad5_ GND EXT2
C6 +5V GND 100n
J5 Net-_J1-Pad3_ GND NC_09 NC_10 Net-_F1-Pad2_ Net-_J1-Pad2_ ESD
.end
