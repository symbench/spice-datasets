.title KiCad schematic
U16 ~RESET NC_01 NC_02 /PCLK NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 /PCLK NC_10 NC_11 ~RESET NC_12 74HC109
U17 ~RESET NC_13 NC_14 /PCLK NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 /PCLK NC_22 NC_23 ~RESET NC_24 74HC109
.end
