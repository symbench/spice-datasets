.title KiCad schematic
J1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 /WAKEA6 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13  
J2 NC_14 NC_15 NC_16 NC_17 /10-INTCCS /SDA /SCL /RX /TX /RESET GND +3V3 VCC +5V  
MODULE1 /TX /RX GND +3V3 +3V3 NC_18 NC_19 NC_20 NC_21 NC_22 GND L80-M39
J4 +3V3 GND /SCL /SDA /WAKEA6 /10-INTCCS /RESET NC_23 CCS811
J3 +3V3 GND /SCL /SDA BME280
.end
