.title KiCad schematic
U2 NC_01 /MotorA/Diagnostic Net-_U2-Pad10_ NC_02 NC_03 Net-_U2-Pad18_ Net-_U2-Pad18_ NC_04 NC_05 Net-_U2-Pad10_ NC_06 /MotorA/Diagnostic NC_07 NC_08 NC_09 NC_10 Net-_U2-Pad17_ Net-_U2-Pad18_ Net-_U2-Pad18_ Net-_U2-Pad17_ NC_11 NC_12 NC_13 NC_14 L6235PD
U3 NC_15 /MotorB/Diagnostic Net-_U3-Pad10_ NC_16 NC_17 Net-_U3-Pad18_ Net-_U3-Pad18_ NC_18 NC_19 Net-_U3-Pad10_ NC_20 /MotorB/Diagnostic NC_21 NC_22 NC_23 NC_24 Net-_U3-Pad17_ Net-_U3-Pad18_ Net-_U3-Pad18_ Net-_U3-Pad17_ NC_25 NC_26 NC_27 NC_28 L6235PD
.end
