.title KiCad schematic
.include "/home/akshay/Downloads/Design_Of_Binary_Phase_Shift_Keying_(bpsk)_Modulator_&_Demodulator_Using_Esim_By_Prof_Raghu_K/Design_Of_BPSK_by_Raghu/BPSK/ZenerD1N750.lib"
V1 ip Net-_R2-Pad2_ sin(0 250)
R1 Net-_C1-Pad1_ ip 470k
C1 Net-_C1-Pad1_ ip 22u
R2 Net-_D2-Pad2_ Net-_R2-Pad2_ 100
C2 GND vd 470u
R3 out vd 100
D5 out GND D1N750
D1 Net-_C1-Pad1_ GND D
D3 vd Net-_C1-Pad1_ D
D4 vd Net-_D2-Pad2_ D
D2 Net-_D2-Pad2_ GND D
.tran .25m 30m
.end
