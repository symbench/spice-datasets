.title KiCad schematic
U$1 /+5V /+5V NC_01 NC_02 NC_03 NC_04 /+5V /+5V /GND NC_05 NC_06 NC_07 /GND /+5V /+5V NC_08 /+12V NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 /+12V /+12V /+12V /GND /GND /GND /GND /GND /GND /GND /GND /GND /GND 581_01_48_005_S
.end
