.title KiCad schematic
P3 GND VCC CONN_VCC
P1 GND GND /BAT /BAT /BAT /BAT /CHARGE /CHARGE GND GND CONN5
U1 GND /BAT VCC TPS61800 module
U2 GND /BAT VCC G5177 module
C1 /BAT GND 47uF
U5 GND /CHG_IN /CHARGE TP5000 Charger
C2 /CHG_IN GND 47uF
U4 GND /BAT VCC LDO_3V5
P2 /CHG_IN /V0.6 /V3.3 NC_01 GND GND USB_Micro
R1 VCC /V3.3 2M
R2 /V3.3 /V0.6 1M
R3 /V0.6 GND 400K
C4 /CHG_IN GND 47uF
P7 /BAT CONN_01X01
P6 GND CONN_01X01
P8 /CHG_IN CONN_01X01
P5 /V0.6 /V3.3 /V3.3 CONN_01X03
P4 /V0.6 /V0.6 /V3.3 CONN_01X03
C3 VCC GND 47uF
C5 /BAT GND 47uF
C6 VCC GND 47uF
.end
