.title KiCad schematic
J2 /Pin1 /Pin2 /Pin3 /Pin4 /Pin5 /Pin6 /Pin7 /Pin8 /Pin9 GND Conn_01x10
J1 /Pin1 /Pin2 /Pin3 /Pin4 /Pin5 /Pin6 /Pin7 /Pin8 /Pin9 Conn_01x09
.end
