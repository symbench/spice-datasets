.title KiCad schematic
D1 5V_L Net-_D1-Pad2_ 5V_L NC_01 WS2812B
D3 5V_L Net-_D3-Pad2_ 5V_L Net-_D1-Pad2_ WS2812B
D5 5V_L Net-_D5-Pad2_ 5V_L Net-_D3-Pad2_ WS2812B
D6 5V_L Net-_D6-Pad2_ 5V_L Net-_D5-Pad2_ WS2812B
D7 5V_L Net-_D7-Pad2_ 5V_L Net-_D6-Pad2_ WS2812B
D8 5V_L Net-_D8-Pad2_ 5V_L Net-_D7-Pad2_ WS2812B
D9 5V_L Net-_D10-Pad4_ 5V_L Net-_D8-Pad2_ WS2812B
D10 5V_L /DOUT..LINK 5V_L Net-_D10-Pad4_ WS2812B
D2 5V_L Net-_D2-Pad2_ GNDL /DOUT..LINK WS2812B
D4 5V_L NC_02 GNDL Net-_D2-Pad2_ WS2812B
C2 GNDL 5V_L C_Small
C4 GNDL 5V_L C_Small
C3 5V_L GNDL C_Small
C1 5V_L 5V_L C_Small
C5 5V_L GNDL C_Small
C6 5V_L GNDL C_Small
C7 5V_L GNDL C_Small
C8 5V_L GNDL C_Small
C9 5V_L GNDL C_Small
C10 5V_L GNDL C_Small
.end
