.title KiCad schematic
U1 Net-_C1-Pad2_ Net-_R1-Pad2_ Net-_R3-Pad2_ 4 Net-_C1-Pad1_ Net-_R4-Pad2_ NC_01 4 LM555
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 0.01u
R1 Net-_J4-Pad1_ Net-_R1-Pad2_ 10k
R5 Net-_R4-Pad2_ Net-_J5-Pad1_ 10k
R4 Net-_C1-Pad2_ Net-_R4-Pad2_ 1M
R2 Net-_R1-Pad2_ Net-_C1-Pad2_ 1M
R3 Net-_Q1-Pad2_ Net-_R3-Pad2_ 10k
R6 Net-_Q1-Pad2_ Net-_C1-Pad2_ 100k
J2 4 Conn_01x01_Male
J3 Net-_J3-Pad1_ Conn_01x01_Male
Q1 Net-_J3-Pad1_ Net-_Q1-Pad2_ Net-_C1-Pad2_ BC547
VCC1 4 Conn_01x01_Male
GND1 Net-_C1-Pad2_ Conn_01x01_Male
J6 4 Conn_01x01_Male
J4 Net-_J4-Pad1_ Conn_01x01_Male
J5 Net-_J5-Pad1_ Conn_01x01_Male
.end
