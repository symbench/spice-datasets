.title KiCad schematic
J1101 +5V +5V +5V +5V /~READ NC_01 /~WRITE /~RESET /A0 /D0 /A1 /D1 /A2 /D2 /A3 /D3 /A4 /D4 /A5 /D5 /A6 /D6 NC_02 /D7 NC_03 Net-_D1101-Pad1_ GNDD GNDD GNDD GNDD GNDD GNDD Conn_02x16_Odd_Even
C1101 GNDD +5V C
C1102 GNDD +5V 100n
D1101 Net-_D1101-Pad1_ /~WAIT D
J1102 +5V +5V +5V +5V /~READ NC_04 /~WRITE /~RESET /A0 /D0 /A1 /D1 /A2 /D2 /A3 /D3 /A4 /D4 /A5 /D5 /A6 /D6 NC_05 /D7 NC_06 Net-_D1102-Pad1_ GNDD GNDD GNDD GNDD GNDD GNDD Conn_02x16_Odd_Even
C1103 GNDD +5V C
C1104 GNDD +5V 100n
D1102 Net-_D1102-Pad1_ /~WAIT D
J1103 +5V +5V +5V +5V /~READ NC_07 /~WRITE /~RESET /A0 /D0 /A1 /D1 /A2 /D2 /A3 /D3 /A4 /D4 /A5 /D5 /A6 /D6 NC_08 /D7 NC_09 Net-_D1103-Pad1_ GNDD GNDD GNDD GNDD GNDD GNDD Conn_02x16_Odd_Even
C1105 GNDD +5V C
C1107 GNDD +5V 100n
D1103 Net-_D1103-Pad1_ /~WAIT D
J1104 +5V +5V +5V +5V /~READ NC_10 /~WRITE /~RESET /A0 /D0 /A1 /D1 /A2 /D2 /A3 /D3 /A4 /D4 /A5 /D5 /A6 /D6 NC_11 /D7 NC_12 Net-_D1104-Pad1_ GNDD GNDD GNDD GNDD GNDD GNDD Conn_02x16_Odd_Even
C1108 GNDD +5V C
C1109 GNDD +5V 100n
D1104 Net-_D1104-Pad1_ /~WAIT D
J1105 +5V +5V +5V +5V /~READ NC_13 /~WRITE /~RESET /A0 /D0 /A1 /D1 /A2 /D2 /A3 /D3 /A4 /D4 /A5 /D5 /A6 /D6 NC_14 /D7 NC_15 Net-_D1105-Pad1_ GNDD GNDD GNDD GNDD GNDD GNDD Conn_02x16_Odd_Even
C1110 GNDD +5V C
C1111 GNDD +5V 100n
D1105 Net-_D1105-Pad1_ /~WAIT D
.end
