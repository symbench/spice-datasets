.title KiCad schematic
J801 GNDD Net-_J801-Pad2_ Net-_J801-Pad3_ Net-_J801-Pad4_ Net-_J801-Pad5_ Net-_J801-Pad6_ FTDI Male
Y801 Net-_C802-Pad1_ Net-_C801-Pad1_ 1.8432MHz
C801 Net-_C801-Pad1_ GNDD 33pF
C802 Net-_C802-Pad1_ GNDD 33pF
C804 GNDD +5V 100nF
C803 GNDD +5V 100pF
U802 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 Net-_C801-Pad1_ GNDD Net-_C802-Pad1_ NC_11 NC_12 NC_13 Net-_U801-Pad3_ NC_14 NC_15 NC_16 NC_17 GNDD Net-_J802-Pad2_ NC_18 Net-_J802-Pad4_ Net-_J802-Pad5_ NC_19 Net-_J802-Pad6_ Net-_U801-Pad10_ +5V +5V NC_20 +5V Net-_U801-Pad2_ NC_21 Net-_J801-Pad2_ NC_22 Net-_J801-Pad5_ Net-_J801-Pad4_ Net-_J801-Pad6_ Net-_U801-Pad4_ +5V +5V +5V ST16C2552_PLCC
R801 Net-_C802-Pad1_ Net-_C801-Pad1_ 680k
U801 Net-_D801-Pad1_ Net-_U801-Pad2_ Net-_U801-Pad3_ Net-_U801-Pad4_ Net-_J801-Pad3_ Net-_J801-Pad3_ Net-_J802-Pad3_ Net-_J802-Pad3_ Net-_U801-Pad10_ 74HC02
D801 Net-_D801-Pad1_ NC_23 D
J802 GNDD Net-_J802-Pad2_ Net-_J802-Pad3_ Net-_J802-Pad4_ Net-_J802-Pad5_ Net-_J802-Pad6_ FTDI Male
R802 GNDD Net-_J801-Pad3_ 4k7
R803 GNDD Net-_J802-Pad3_ 4k7
.end
