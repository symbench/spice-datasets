.title KiCad schematic
IC1 Net-_C5-Pad2_ Net-_C1-Pad1_ Net-_IC1-Pad3_ Net-_IC1-Pad4_ /FB Net-_C7-Pad1_ GND Net-_C5-Pad1_ GND TPS54560BDDAR
R2 Net-_IC1-Pad3_ GND 80.6k
R1 Net-_C1-Pad1_ Net-_IC1-Pad3_ 1050k
C4 Net-_C1-Pad1_ GND 1210B225K101CT
C3 Net-_C1-Pad1_ GND 1210B225K101CT
C2 Net-_C1-Pad1_ GND 1210B225K101CT
C1 Net-_C1-Pad1_ GND 1210B225K101CT
C8 /12V+ GND EMK325BJ226KM-P
C9 /12V+ GND EMK325BJ226KM-P
C10 /12V+ GND EMK325BJ226KM-P
L1 Net-_C5-Pad1_ /12V+ PA4343.133NLT
D1 Net-_C5-Pad1_ GND B560C-13-F
R4 Net-_C7-Pad1_ Net-_C6-Pad1_ 13k
C6 Net-_C6-Pad1_ GND 4700pF
R5 /12V+ /FB 143k
R6 /FB GND 10.2k
C7 Net-_C7-Pad1_ GND 47pF
C5 Net-_C5-Pad1_ Net-_C5-Pad2_ 100nF_min8V
R3 Net-_IC1-Pad4_ GND 162k
.end
