.title KiCad schematic
U201 COM COM COM COM COM COM COM COM COM COM COM COM COM COM COM COM COM COM PP_VDD_SOC_CAP PP_VDD_ARM_CAP PP_VDD_ARM_CAP PP_VDD_ARM_CAP COM COM COM PP_VDD_SOC_CAP PP_VDD_SOC_IN PP_VDD_SOC_IN PP_VDD_ARM_CAP COM COM COM PP_VDD_SOC_CAP PP_VDD_SOC_IN PP_VDD_SOC_IN PP_VDD_SOC_CAP COM COM PP_VDD_SOC_CAP PP_VDD_SOC_IN PP_VDD_SOC_IN PP_VDD_SOC_CAP COM COM COM PP_VDD_SOC_CAP PP_VDD_SOC_CAP PP_VDD_SOC_CAP PP_VDD_SOC_CAP COM PP_VDDA_ADC_3P3 COM COM COM COM COM COM PP_VDDA_ADC_3P3 COM COM PP_VDD_SNVS_CAP PP_VDD_HIGH_IN PP_VDD_SNVS_IN PP_NVCC_PLL COM COM COM COM PP_VDD_HIGH_CAP PP_VDD_HIGH_CAP COM COM COM COM COM COM MCIMX6Y2DVM
C208 PP_VDD_SOC_IN COM 0.22u
C211 PP_VDD_SOC_IN COM 22u
C209 PP_VDD_SOC_IN COM 0.22u
C210 PP_VDD_SOC_IN COM 10u
C201 PP_VDD_ARM_CAP COM 0.22u
C202 PP_VDD_ARM_CAP COM 0.22u
C203 PP_VDD_ARM_CAP COM 22u
C204 PP_VDD_SOC_CAP COM 0.22u
C205 PP_VDD_SOC_CAP COM 0.22u
C207 PP_VDD_SOC_CAP COM 22u
C206 PP_VDD_SOC_CAP COM 0.22u
C212 PP_VDD_HIGH_IN COM 0.22u
C213 PP_VDD_HIGH_IN COM 10u
C214 PP_VDD_HIGH_CAP COM 0.22u
C215 PP_VDD_HIGH_CAP COM 10u
C218 PP_VDD_SNVS_IN COM 0.22u
C219 PP_VDD_SNVS_CAP COM 0.22u
C216 PP_NVCC_PLL COM 0.22u
C217 PP_NVCC_PLL COM 10u
.end
