.title KiCad schematic
U1 /RST /RXD /TXD /ZERO_CROSS /TRIAC_GATE /LED_RUNNING +5V GND Net-_C3-Pad2_ Net-_C4-Pad1_ /FAN_S /CLK /CS /SO /SW_STOP_MODE /SW_START_SET /MOSI /MISO /SCK +5V +5V GND /A0 /A1 NC_01 NC_02 /SDA /SCL ATmega328P-PU
Y1 Net-_C3-Pad2_ Net-_C4-Pad1_ 16MHz
C3 GND Net-_C3-Pad2_ 22p
C4 Net-_C4-Pad1_ GND 22p
J1 +5V GND PWR_IN
C2 GND +5V 15p
C1 GND +5V 15p
R2 +5V /RST 4k7
D2 +5V /RST 5.1V
C5 GND /RST 15p
R3 Net-_R3-Pad1_ /RST 330
SW1 Net-_R3-Pad1_ GND SW_RST
J2 /MOSI +5V NC_03 GND /RST GND /SCK GND /MISO GND SPI
R1 Net-_D1-Pad1_ GND 1k
D1 Net-_D1-Pad1_ +5V PWR
J3 /SDA /SCL GND +5V DISP
J5 GND +5V /CLK /CS /SO THERM
J6 +5V GND /FAN_S FAN
J7 +5V GND /ZERO_CROSS /TRIAC_GATE HEAT
J4 +5V GND /RXD /TXD UART
RV1 +5V /A0 GND 100K_VAL
RV2 +5V /A1 GND 100K_PAR
SW2 /SW_STOP_MODE GND SW_STOP_MODE
SW3 /SW_START_SET GND SW_START_SET
R4 Net-_D3-Pad1_ GND 1k
D3 Net-_D3-Pad1_ /LED_RUNNING RUN
.end
