.title KiCad schematic
U15 NC_01 NC_02 Net-_U15-Pad3_ NC_03 NC_04 NC_05 NC_06 Net-_U15-Pad3_ NC_07 NC_08 SC39-11
U17 NC_09 NC_10 Net-_U17-Pad3_ NC_11 NC_12 NC_13 NC_14 Net-_U17-Pad3_ NC_15 NC_16 SC39-11
U19 NC_17 NC_18 Net-_U19-Pad3_ NC_19 NC_20 NC_21 NC_22 Net-_U19-Pad3_ NC_23 NC_24 SC39-11
U21 NC_25 NC_26 Net-_U21-Pad3_ NC_27 NC_28 NC_29 NC_30 Net-_U21-Pad3_ NC_31 NC_32 SC39-11
U23 NC_33 NC_34 Net-_U23-Pad3_ NC_35 NC_36 NC_37 NC_38 Net-_U23-Pad3_ NC_39 NC_40 SC39-11
U25 NC_41 NC_42 Net-_U25-Pad3_ NC_43 NC_44 NC_45 NC_46 Net-_U25-Pad3_ NC_47 NC_48 SC39-11
CN1 NC_49 NC_50 NC_51 NC_52 NC_53 NC_54 NC_55 NC_56 NC_57 0.1µF
CN2 NC_58 NC_59 NC_60 NC_61 NC_62 NC_63 NC_64 NC_65 NC_66 0.1µF
CN3 NC_67 NC_68 NC_69 NC_70 NC_71 NC_72 NC_73 NC_74 NC_75 0.1µF
.end
