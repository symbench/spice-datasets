.title KiCad schematic
J1 GND +12V_BUS NC_01 Net-_J1-Pad4_ Conn_01x04
Q1 /PWM_01 GND Net-_J1-Pad4_ 2N7002
R6 /PWM_01 GND 10K
R1 +5V_BUS Net-_J1-Pad4_ 4.7K
J2 GND +12V_BUS NC_02 Net-_J2-Pad4_ Conn_01x04
Q2 /PWM_02 GND Net-_J2-Pad4_ 2N7002
R7 /PWM_02 GND 10K
R2 +5V_BUS Net-_J2-Pad4_ 4.7K
J3 GND +12V_BUS NC_03 Net-_J3-Pad4_ Conn_01x04
Q3 /PWM_03 GND Net-_J3-Pad4_ 2N7002
R8 /PWM_03 GND 10K
R3 +5V_BUS Net-_J3-Pad4_ 4.7K
J4 GND +12V_BUS NC_04 Net-_J4-Pad4_ Conn_01x04
Q4 /PWM_04 GND Net-_J4-Pad4_ 2N7002
R9 /PWM_04 GND 10K
R4 +5V_BUS Net-_J4-Pad4_ 4.7K
J5 GND +12V_BUS NC_05 Net-_J5-Pad4_ Conn_01x04
Q5 /PWM_05 GND Net-_J5-Pad4_ 2N7002
R10 /PWM_05 GND 10K
R5 +5V_BUS Net-_J5-Pad4_ 4.7K
C4 +12V_BUS GND 100uF
C2 +12V_BUS GND 100uF
C3 +5V_BUS GND 100pF
C5 +5V_BUS GND 100uF
C1 +12V_BUS GND 100pF
.end
