.title KiCad schematic
J49 GND /SDIO_DATA_0 /SDIO_DATA_CLK /SDIO_DATA_1 GND /SDIO_DATA_2 /SDIO_DATA_CMD /SDIO_DATA_3 /WL_REG_ON /CLK32K /WL_WAKE_AP GND /VCC /VCC SBBJ49
J50 NC_01 /BT_UART_RX NC_02 /BT_UART_TX NC_03 /BT_UART_CTS NC_04 /BT_UART_RTS GND GND /BT_WAKE_AP /BT_RST_N /AP_WAKE_BT /VDDIO GND GND SBBJ50
U1 GND Net-_J1-Pad1_ GND GND GND GND GND GND Net-_J2-Pad1_ GND GND NC_05 Net-_C2-Pad1_ Net-_C1-Pad1_ /WL_REG_ON /WL_WAKE_AP /SDIO_DATA_CMD /SDIO_DATA_CLK /SDIO_DATA_3 /SDIO_DATA_2 /SDIO_DATA_0 /SDIO_DATA_1 GND Net-_R1-Pad2_ Net-_C3-Pad1_ Net-_L1-Pad1_ NC_06 NC_07 NC_08 NC_09 /CLK32K GND NC_10 /VDDIO NC_11 /VCC NC_12 /BT_RST_N GND /BT_UART_TX /BT_UART_RX /BT_UART_RTS /BT_UART_CTS NC_13 NC_14 NC_15 NC_16 NC_17 /AP_WAKE_BT /BT_WAKE_AP ap6356s
Y1 Net-_C1-Pad1_ GND Net-_C2-Pad1_ GND 37.4MHz, 1.6x1.2mm, Epson FA-118T
C1 Net-_C1-Pad1_ GND C
C2 Net-_C2-Pad1_ GND C
J1 Net-_J1-Pad1_ GND GND UFL
J2 Net-_J2-Pad1_ GND GND UFL
C3 Net-_C3-Pad1_ GND 4.7u, 0603, X5R, 10V
R1 /VDDIO Net-_R1-Pad2_ 10K, 1%
L1 Net-_L1-Pad1_ Net-_C3-Pad1_ 4.7uH, 1A
C4 /VCC GND 1uF
C5 /VCC GND 4.7uF
.end
