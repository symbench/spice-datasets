.title KiCad schematic
U1 NC_01 NC_02 Net-_U1-Pad3_ NC_03 NC_04 NC_05 NC_06 Net-_U1-Pad3_ NC_07 NC_08 SC39-11
.end
