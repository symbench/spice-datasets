.title KiCad schematic
U1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 /~reset NC_07 NC_08 NC_09 NC_10 GND +3V3 NC_11 NC_12 NC_13 NC_14 GND +3V3 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 GND +3V3 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 /swdio GND +3V3 /swdclk NC_39 NC_40 NC_41 NC_42 NC_43 NC_44 NC_45 NC_46 NC_47 NC_48 NC_49 NC_50 NC_51 GND +3V3 STM32F091RCTx
C9 /~reset GND 100n
C1 +3V3 GND 100n
C2 +3V3 GND 100n
C3 +3V3 GND 100n
C4 +3V3 GND 100n
C5 +3V3 GND 10n
C6 +3V3 GND 4.7u
C7 +3V3 GND 4.7u
C8 +3V3 GND 1u
J1 +3V3 /swdio GND /swdclk GND NC_52 NC_53 NC_54 GND /~reset ARM_JTAG_SWD_10
.end
