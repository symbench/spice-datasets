.title KiCad schematic
M1 NC_01 NC_02 DriveMotor
.end
