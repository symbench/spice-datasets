.title KiCad schematic
U1 +5V GNDREF NC_01 NC_02 GNDREF ACS754
.end
