.title KiCad schematic
J4 GND +3V3 CS_3V3 CLK_3V3 MISO_3V3 MOSI_3V3 IN
U3 GND +1V8 +3V3 AP1117-18
C2 +1V8 GND 100nF
C1 +3V3 GND 100nF
U1 GND +1V8 MOSI_1V8 MISO_1V8 MISO_3V3 MOSI_3V3 Net-_C3-Pad1_ Net-_C3-Pad1_ GTL2002DP
U2 GND +1V8 CLK_1V8 CS_1V8 CS_3V3 CLK_3V3 Net-_C4-Pad1_ Net-_C4-Pad1_ GTL2002DP
J3 MOSI_1V8 MISO_1V8 CLK_1V8 CS_1V8 +1V8 GND OUT
R3 MOSI_1V8 +1V8 3K3
R1 MISO_1V8 +1V8 3K3
R4 CLK_1V8 +1V8 3K3
R2 CS_1V8 +1V8 3K3
R7 MOSI_3V3 +3V3 3K3
R9 MISO_3V3 +3V3 3K3
R8 CLK_3V3 +3V3 3K3
R5 CS_3V3 +3V3 3K3
C3 Net-_C3-Pad1_ GND 100nF
C4 Net-_C4-Pad1_ GND 100nF
R6 Net-_C4-Pad1_ +3V3 200K
R10 Net-_C3-Pad1_ +3V3 200K
R11 Net-_D1-Pad2_ +3V3 3K3
D1 GND Net-_D1-Pad2_ LED
J1 GND +1V8 +1V8 +1V8 GND GND PWR
.end
