.title KiCad schematic
Y1 NC_01 NC_02 Crystal
U1 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 GND NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 GND NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 GND NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 GND NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 GND NC_43 GND NC_44 FT2232D
.end
