.title KiCad schematic
BT1 Net-_BT1-Pad1_ Net-_BT1-Pad2_ Battery_Cell
R1 Net-_BT1-Pad1_ Net-_BT1-Pad2_ R
.end
