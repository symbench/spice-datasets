.title KiCad schematic
U3 NC_01 COM_DATA GND CH1_DATA 3.3V 74LVC1G125
U4 NC_02 CH1_DATA GND COM_DATA 3.3V 74LVC1G125
U5 NC_03 COM_DATA GND CH2_DATA 3.3V 74LVC1G125
U6 NC_04 CH2_DATA GND COM_DATA 3.3V 74LVC1G125
U7 NC_05 COM_DATA GND CH3_DATA 3.3V 74LVC1G125
U8 NC_06 CH3_DATA GND COM_DATA 3.3V 74LVC1G125
.end
