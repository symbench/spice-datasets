.title KiCad schematic
J2 GND GND +5V +5V GND +3V3 +3V3 GND GP21 GP20 SD_D2 GND GP19 GP16 GP13 GND GP12 GP6 GP5 GND ID_SC ID_SD SCK GND CS0 CS1 MISO MOSI GND SD_D1 SD_D0 GND SD_CLK SD_CMD SD_D3 GND GP18 RX TX GND GP17 GP4 SCL SDA GND +3V3 +3V3 GND +5V +5V GND Conn_01x50_shd
J1 +3V3 +5V SDA +5V SCL GND GP4 TX GND RX GP17 GP18 SD_D3 GND SD_CLK SD_CMD +3V3 SD_D0 MOSI GND MISO SD_D1 SCK CS0 GND CS1 ID_SD ID_SC GP5 GND GP6 GP12 GP13 GND GP19 GP16 SD_D2 GP20 GND GP21 RPi
J3 GND GND +5V +5V GND +3V3 +3V3 GND GP21 GP20 SD_D2 GND GP19 GP16 GP13 GND GP12 GP6 GP5 GND ID_SC ID_SD SCK GND CS0 CS1 MISO MOSI GND SD_D1 SD_D0 GND SD_CLK SD_CMD SD_D3 GND GP18 RX TX GND GP17 GP4 SCL SDA GND +3V3 +3V3 GND +5V +5V GND Conn_01x50_shd
.end
