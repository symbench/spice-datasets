.title KiCad schematic
U3 /Coil /Coil_Out +BATT NC_01 /Power_Out V23074A2002A403
U2 /Coil /Coil_Out +BATT NC_02 /Fun_Out V23074A2002A403
P6 GNDPWR +BATT POWER_IN
R7 +BATT Net-_D2-Pad1_ 4.7k
R8 /24v Net-_D3-Pad1_ 4.7k
D2 Net-_D2-Pad1_ GNDPWR LED
D3 Net-_D3-Pad1_ GNDPWR LED
R9 +12V Net-_D4-Pad1_ 2.2k
D4 Net-_D4-Pad1_ GND LED
D5 Net-_D5-Pad1_ GNDPWR LED
R10 /Coil Net-_D5-Pad1_ 4.7k
U1 GNDPWR GNDPWR /24v GND NC_03 +12V CCG30-24-xxS
C3 GNDPWR /24v 470
C6 +12V GND 470
P4 GND +12V 12v
C1 +12V GND 0.1u
P5 GND +12V 12v
C2 +12V GND 0.1u
P3 Net-_D1-Pad2_ /24v POW_SW
P7 GNDPWR FRAMEGND
IC1 Net-_IC1-Pad1_ GND Net-_IC1-Pad3_ Net-_IC1-Pad4_ TLP291
IC2 Net-_IC2-Pad1_ GNDPWR GND /Relay_state TLP291
R1 /24v Net-_IC1-Pad4_ 2.2k
R2 Net-_IC2-Pad1_ /Coil 4.7k
P8 GND +12V /Forced_shutdown /Relay_state main-signal
C4 GND +12V 0.1u
R6 +12V /Relay_state 10k
R5 /Relay_state GND 2.2k
R4 /Forced_shutdown Net-_IC1-Pad1_ 330
R3 Net-_IC1-Pad3_ GNDPWR 2.2k
Q1 Net-_IC1-Pad3_ GNDPWR /Coil_Out MOSFET_N_123
JP1 GNDPWR /Coil_Out JUMPER
P2 /Coil Net-_P1-Pad1_ EMERGENCY
P1 Net-_P1-Pad1_ /24v EMERGENCY
P10 GNDPWR /Power_Out POWER_OUT
P11 GNDPWR /Fun_Out FUN_OUT
P9 GND +12V /Forced_shutdown /Relay_state main-signal
C5 GND +12V 0.1u
D6 Net-_D6-Pad1_ GNDPWR LED
R11 /Power_Out Net-_D6-Pad1_ 4.7k
D7 Net-_D7-Pad1_ GNDPWR LED
R12 /Fun_Out Net-_D7-Pad1_ 4.7k
D1 +BATT Net-_D1-Pad2_ DIODE
.end
