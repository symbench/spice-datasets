.title KiCad schematic
U1 GND +3V3 EN NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 GND NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 GPIO0 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 SCL RX TX SDA NC_28 GND GND ESP32-WROVER
Q2 Net-_Q2-Pad1_ /DTR GPIO0 BC847
Q1 Net-_Q1-Pad1_ /CTS EN BC847
R1 /DTR Net-_Q1-Pad1_ 10K
R2 /CTS Net-_Q2-Pad1_ 10K
J1 GND /CTS +3V3 RX TX /DTR PROGRAMMING
C4 +3V3 GND 100pF
C1 +3V3 GND 10uF
C2 +3V3 GND 10uF
C3 +3V3 GND 100pF
R3 +3V3 SDA 4K7
R4 +3V3 SCL 4k7
J2 NC_29 +5V GND TX RX GND MainIO
.end
