.title KiCad schematic
U1 NC_01 +5V NC_02 GND NC_03 AD8331EVALZ
.end
