.title KiCad schematic
P1 3.3V 5v NC_01 5v NC_02 GND NC_03 NC_04 GND NC_05 NC_06 NC_07 NC_08 GND NC_09 NC_10 3.3V NC_11 NC_12 GND NC_13 NC_14 NC_15 NC_16 GND NC_17 NC_18 NC_19 GPIO05 GND GPIO06 DIR_1 NC_20 GND NC_21 GPIO16 NC_22 DIR_2 GND GPIO21 Raspberry Pi Zero W
P2 GND DIR_1 5v GPIO16 1B_1 Net-_P2-Pad6_ 1A_1 Net-_P2-Pad6_ 2A_1 NC_23 2B_1 NC_24 GND NC_25 Battery+ GPIO05 STEPPER_1
C1 Battery+ GND 470uF
P4 2B_1 2A_1 1A_1 1B_1 MOTOR 1
P3 GND DIR_2 5v GPIO21 1B_2 Net-_P3-Pad6_ 1A_2 Net-_P3-Pad6_ 2A_2 NC_26 2B_2 NC_27 GND NC_28 Battery+ GPIO06 STEPPER_2
C2 Battery+ GND 470uF
P5 2B_2 2A_2 1A_2 1B_2 MOTOR 2
P6 Battery+ Battery- PWR
D1 Net-_D1-Pad1_ 5v LED
R1 Net-_D1-Pad1_ GND 330
U1 Battery+ Battery+ Battery- Battery- Net-_SW1-Pad2_ Net-_SW1-Pad2_ GND GND LM2596_mini_module
SW1 NC_29 Net-_SW1-Pad2_ 5v Switch_SPDT_x2
.end
