.title KiCad schematic
J1 GND +BATT Net-_J1-Pad3_ Net-_J1-Pad3_ Conn_02x02_Counter_Clockwise
U2 GND +3V3 +BATT AZ1117-3.3
U3 GND +5V +BATT AZ1117-5.0
U4 GND +5V +BATT AZ1117-5.0
U1 GND +3V3 +BATT AZ1117-3.3
J2 NC_01 +5V +3V3 GND Conn_01x04_Female
J3 NC_02 +5V +3V3 GND Conn_01x04_Female
J4 NC_03 +5V +3V3 GND Conn_01x04_Female
J5 NC_04 +5V +3V3 GND Conn_01x04_Female
J6 NC_05 +5V +3V3 GND Conn_01x04_Female
C1 +BATT GND CAP
C2 +3V3 GND CAP
C3 +5V GND CAP
R1 +BATT Net-_D1-Pad1_ R
D1 Net-_D1-Pad1_ GND LED
C4 +3V3 GND CAP
C5 +5V GND CAP
C6 +BATT GND CAP
C7 +BATT GND CAP
C8 +BATT GND CAP
.end
