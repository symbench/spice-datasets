.title KiCad schematic
U1 Net-_C2-Pad1_ Net-_R1-Pad1_ Net-_R1-Pad1_ Net-_J1-Pad24_ GND NC_01 GND NC_02 GND NC_03 GND NC_04 GND VCC 74HC14
R1 Net-_R1-Pad1_ Net-_C2-Pad1_ 1M
R2 Net-_C1-Pad1_ Net-_R1-Pad1_ 10k
Y1 Net-_C2-Pad1_ Net-_C1-Pad1_ 4MHz Crystal
C1 Net-_C1-Pad1_ GND 3.3p
C2 Net-_C2-Pad1_ GND 3.3p
C3 VCC GND 0.1u
J1 VCC NC_05 GND NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 GND NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 GND Net-_J1-Pad24_ Conn_01x24_Female
.end
