.title KiCad schematic
BATT1 VLIPO GND JST 2PH
X2 /CC1 /D+ /D- NC_01 GND /VUSB /CC2 /D+ /D- NC_02 GND /VUSB USB Type C
D2 /VUSB VBUS SK34A
R1 GND /CC2 5.1K
R2 GND /CC1 5.1K
D4 /OUT Net-_D4-PadC_ RED
R7 /CHG Net-_D4-PadC_ 10K
C7 VLIPO GND 10uF
C2 VBUS GND 10uF
C4 /OUT GND 10uF
C5 /OUT GND 10uF
U$1 MOUNTINGHOLE2.5
U$3 MOUNTINGHOLE2.5
U$2 MOUNTINGHOLE2.5
U$4 MOUNTINGHOLE2.5
X1 Net-_D1-PadA_ Net-_D1-PadA_ GND GND 2.1mm DC
SYSOUT1 /OUT GND JST 2PH
D1 Net-_D1-PadA_ VBUS SK34A
R3 /ISET Net-_1.5A1-Pad2_ 590
C1 VBUS GND 10uF
R5 /ISET Net-_0.5A1-Pad2_ 2K
1.5A1 GND Net-_1.5A1-Pad2_ SOLDERJUMPER
0.5A1 GND Net-_0.5A1-Pad2_ SOLDERJUMPER
R4 /ISET Net-_1A1-Pad2_ 1K
1A1 GND Net-_1A1-Pad2_ SOLDERJUMPERCLOSED
X3 /THERM VLIPO VLIPO /CE /EN2 /EN1 /PGOOD GND /CHG /OUT /OUT /ILIM VBUS GND /ITERM /ISET GND BQ24074
D3 /OUT Net-_D3-PadC_ GREEN
R8 /ILIM GND 1K
R9 /ITERM GND 10K
JP2 GND VLIPO GND /OUT /CHG /PGOOD /CE /ISET /THERM GND VBUS HEADER-1X1176MIL
C3 /OUT GND 10uF
C6 VLIPO GND 10uF
JP1 /D+ /D- HEADER-1X2ROUND
FID3 FIDUCIAL_1MM
FID2 FIDUCIAL_1MM
FID1 FIDUCIAL_1MM
R11 Net-_R11-Pad1_ GND 10K
SJ2 /OUT /EN2 GND SOLDERJUMPER_2WAY
SJ1 /OUT /EN1 GND SOLDERJUMPER_2WAY
R6 /PGOOD Net-_D3-PadC_ 10K
R10 /CE GND 10K
THERM1 Net-_R11-Pad1_ /THERM SOLDERJUMPERCLOSED
JP4 GND HEADER-1X1
JP3 VBUS HEADER-1X1
.end
