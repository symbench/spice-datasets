.title KiCad schematic
J3 NC_01 /P5V_HAT NC_02 /P5V_HAT NC_03 /GND NC_04 NC_05 /GND NC_06 NC_07 NC_08 NC_09 /GND NC_10 NC_11 NC_12 NC_13 NC_14 /GND NC_15 NC_16 NC_17 NC_18 /GND NC_19 /ID_SD_EEPROM /ID_SC_EEPROM NC_20 /GND NC_21 NC_22 NC_23 /GND NC_24 NC_25 NC_26 NC_27 /GND NC_28 40HAT
Q1 Net-_Q1-Pad1_ /P5V_HAT /P5V DMG2305UX
Q2 Net-_Q2-Pad1_ Net-_Q2-Pad1_ Net-_Q2-Pad1_ Net-_Q1-Pad1_ /P5V_HAT /P5V DMMT5401
U2 Net-_U2-Pad1_ Net-_U2-Pad1_ Net-_U2-Pad1_ NC_29 /ID_SD_EEPROM /ID_SC_EEPROM NC_30 NC_31 CAT24C32
.end
