.title KiCad schematic
U1 GND +3V3 +5V +3V3 LM1117-3.3
C2 +3V3 GND CP
C3 +3V3 GND C
CON1 +5V GND MISO MOSI RXD SCK SCL SDA SSEL TXD UEXT-5V
J1 +3V3 +5V GND TXD RXD SCL SDA MISO MOSI SCK SSEL CONN_01X11
C1 +5V GND CP
.end
