.title KiCad schematic
U2 SCL SDA NC_01 3.3V GND NRST NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 Net-_U1-Pad4_ NC_10 NC_11 NC_12 NC_13 NC_14 STM32G030F6P6
R3 3.3V NRST R_US
SW1 GND NRST SW_Push
R1 3.3V SCL R_US
R2 3.3V SDA R_US
U1 5V GND NC_15 Net-_U1-Pad4_ GND 3.3V SN74LVC1T45DBVR
.end
