.title KiCad schematic
U1 BASE EMITTER COLLECTOR MJD210
P1 COLLECTOR EMITTER BASE CONN_01X03
.end
