.title KiCad schematic
C98 NC_01 Net-_C100-Pad2_ C
C100 NC_02 Net-_C100-Pad2_ C
C99 Net-_C101-Pad1_ NC_03 C
C101 Net-_C101-Pad1_ NC_04 C
J36 Net-_C100-Pad2_ NC_05 Net-_C102-Pad2_ Net-_C103-Pad2_ NC_06 Net-_C101-Pad1_ InConnector
J37 Net-_C106-Pad2_ NC_07 Net-_C104-Pad1_ Net-_C105-Pad1_ NC_08 Net-_C107-Pad1_ OutConnector
U21 NC_09 Net-_R244-Pad1_ Net-_C102-Pad1_ NC_10 NC_11 Net-_C104-Pad2_ NC_12 NC_13 OPA333xxD
R248 NC_14 Net-_C102-Pad1_ R
R246 Net-_C102-Pad2_ Net-_C104-Pad1_ R
R244 Net-_R244-Pad1_ Net-_C102-Pad2_ R
C104 Net-_C104-Pad1_ Net-_C104-Pad2_ C
C102 Net-_C102-Pad1_ Net-_C102-Pad2_ C
R250 Net-_R244-Pad1_ Net-_C104-Pad2_ R
U22 NC_15 Net-_R245-Pad1_ Net-_C103-Pad1_ NC_16 NC_17 Net-_C105-Pad2_ NC_18 NC_19 OPA333xxD
R249 NC_20 Net-_C103-Pad1_ R
R247 Net-_C103-Pad2_ Net-_C105-Pad1_ R
R245 Net-_R245-Pad1_ Net-_C103-Pad2_ R
C105 Net-_C105-Pad1_ Net-_C105-Pad2_ C
C103 Net-_C103-Pad1_ Net-_C103-Pad2_ C
R251 Net-_R245-Pad1_ Net-_C105-Pad2_ R
C106 NC_21 Net-_C106-Pad2_ C
C108 NC_22 Net-_C106-Pad2_ C
C107 Net-_C107-Pad1_ NC_23 C
C109 Net-_C107-Pad1_ NC_24 C
.end
