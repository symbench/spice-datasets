.title KiCad schematic
C2 +3V3 GND 0.1u
U1 GND GND GND GND /SDA /SCL GND +3V3 CK_CUSTOM_M24M02-DRMN6TP
R3 +3V3 /SCL 4.7k
R4 +3V3 /SDA 4.7k
R2 /SDA +3V3 4.7k
R1 /SCL +3V3 4.7k
C1 +3V3 NC_01 0.1u
.end
