.title KiCad schematic
U1 Net-_R5-Pad2_ rtcVcc gnd vcc gnd vcc NC_01 NC_02 NC_03 NC_04 busy reset d.c cs d11 d12 d13 vcc NC_05 vcc gnd NC_06 NC_07 NC_08 NC_09 NC_10 sda scl d10 NC_11 NC_12 NC_13 ATMEGA328P-AU
R1 d10 vcc R
SW1 Net-_R5-Pad2_ vcc Switch_SW_Push
R5 gnd Net-_R5-Pad2_ R
IC1 NC_14 rtcVcc NC_15 gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd Net-_BT2-Pad1_ sda scl DS3231
R2 rtcVcc gnd R
R3 vcc scl R
R4 vcc sda R
L1 vcc Net-_C3-Pad2_ INDUCTOR
C2 vcc gnd C
Q1 gdr rese Net-_C3-Pad2_ 2N7000 switched S and G due to footprint
C3 Net-_C3-Pad1_ Net-_C3-Pad2_ C
D3 prevgh Net-_C3-Pad2_ MBR0530
D2 Net-_C3-Pad1_ prevgl MBR0530
D1 gnd Net-_C3-Pad1_ MBR0530
R6 gdr gnd R
R7 rese gnd R
J2 NC_16 gdr rese Net-_C13-Pad1_ Net-_C12-Pad1_ NC_17 NC_18 gnd busy reset d.c cs d13 d11 vcc vcc gnd Net-_C8-Pad1_ Net-_C5-Pad1_ Net-_C9-Pad1_ prevgh Net-_C10-Pad1_ prevgl Net-_C11-Pad1_ otp_FPC24
C13 Net-_C13-Pad1_ gnd C
C12 Net-_C12-Pad1_ gnd C
C8 Net-_C8-Pad1_ gnd C
C5 Net-_C5-Pad1_ gnd C
C9 Net-_C9-Pad1_ gnd C
C6 prevgh gnd C
C10 Net-_C10-Pad1_ gnd C
C7 prevgl gnd C
C11 Net-_C11-Pad1_ gnd C
C4 vcc gnd C
J1 d13 d12 d11 d10 gnd vcc Conn_01x06_Female
BT1 vcc gnd Battery_Cell
C1 vcc gnd C
BT2 Net-_BT2-Pad1_ gnd Battery_Cell
.end
