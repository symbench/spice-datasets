.title KiCad schematic
U3 /NX2_8 /NX2_9 /A2 /D2 +5V /B2 /C2 /NX2_2 /NX2_3 /NX2_7 /NX2_6 GND /NX2_4 /NX2_5 /NX2_1 /NX2_0 74141
U1 /B1 /C1 /D1 /A2 /B2 /C2 /D2 GND /SEROUT +5V /CLK /LATCH /nOE /DATA /A1 +5V 74HC595
NX2 /NX2_0 /NX2_1 /NX2_2 /NX2_3 /NX2_4 /NX2_5 /NX2_6 /NX2_7 /NX2_8 /NX2_9 /NX2_Anode IN-12A
R2 /NX2_Anode /+170V 12k
NX1 /NX1_0 /NX1_1 /NX1_2 /NX1_3 /NX1_4 /NX1_5 /NX1_6 /NX1_7 /NX1_8 /NX1_9 /NX1_Anode IN-12A
R1 /NX1_Anode /+170V 12k
J1 +5V GND /SEROUT NC_01 /+170V /nOE /DATA /CLK /LATCH Conn_01x09_Male
U2 /NX1_8 /NX1_9 /A1 /D1 +5V /B1 /C1 /NX1_2 /NX1_3 /NX1_7 /NX1_6 GND /NX1_4 /NX1_5 /NX1_1 /NX1_0 74141
.end
