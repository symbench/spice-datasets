.title KiCad schematic
U1 /A0 /A1 /A2 /O0 /O1 /O2 /O3 GND /O4 /O5 /O6 /O7 INT SCL SDA VCC PCF8574
J1 VCC SDA SCL INT GND I2C
C1 VCC GND 100nF
D1 /O0 Net-_D1-Pad2_ LED
R2 VCC Net-_D1-Pad2_ 1K
D2 /O1 Net-_D2-Pad2_ LED
R3 VCC Net-_D2-Pad2_ 1K
D3 /O2 Net-_D3-Pad2_ LED
R4 VCC Net-_D3-Pad2_ 1K
D4 /O3 Net-_D4-Pad2_ LED
R5 VCC Net-_D4-Pad2_ 1K
D5 /O4 Net-_D5-Pad2_ LED
R6 VCC Net-_D5-Pad2_ 1K
D6 /O5 Net-_D6-Pad2_ LED
R7 VCC Net-_D6-Pad2_ 1K
D7 /O6 Net-_D7-Pad2_ LED
R8 VCC Net-_D7-Pad2_ 1K
D8 /O7 Net-_D8-Pad2_ LED
R9 VCC Net-_D8-Pad2_ 1K
JP3 VCC /A2 GND A0
JP2 VCC /A1 GND A1
JP1 VCC /A0 GND A2
J2 VCC /O0 /O1 /O2 /O3 /O4 /O5 /O6 /O7 GND IO
R1 VCC INT 10K
R10 VCC SDA 10K
R11 VCC SCL 10K
.end
