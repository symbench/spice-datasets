.title KiCad schematic
J1 GND 3V3 EN SENSOR_VP SENSOR_VN IO34 IO35 IO32 IO33 IO25 IO26 IO27 IO14 IO12 IO13 SD2 SD3 CMD Conn_01x18
J2 GND IO23 IO22 TXD0 RXD0 IO21 IO19 IO18 IO5 IO17 IO16 IO4 IO0 IO2 IO15 SD1 SD0 CLK Conn_01x18
U1 GND 3V3 EN SENSOR_VP SENSOR_VN IO34 IO35 IO32 IO33 IO25 IO26 IO27 IO14 IO12 GND IO13 SD2 SD3 CMD CLK SD0 SD1 IO15 IO2 IO0 IO4 IO16 IO17 IO5 IO18 IO19 GND IO21 RXD0 TXD0 IO22 IO23 GND GND ESP32-WROOM-32
C1 3V3 GND 22uF
C2 3V3 GND 22uF
SW1 GND EN SW_Push
C3 EN GND 0.1uF
SW2 GND IO0 SW_Push
C4 IO0 GND 0.1uF
.end
