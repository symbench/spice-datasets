.title KiCad schematic
N2 V20190807
N1 OHWLOGO
U1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 LT1021__H
.end
