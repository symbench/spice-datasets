.title KiCad schematic
U7 NC_01 NC_02 NC_03 Net-_U6-Pad4_ Net-_U6-Pad6_ NC_04 Net-_U6-Pad5_ Net-_U6-Pad18_ NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 Net-_U6-Pad21_ Net-_U6-Pad17_ NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 Net-_U6-Pad19_ NC_27 NC_28 NC_29 NC_30 Net-_U6-Pad22_ NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 SC16C2550BIB48
U6 NC_41 NC_42 NC_43 Net-_U6-Pad4_ Net-_U6-Pad5_ Net-_U6-Pad6_ NC_44 NC_45 NC_46 NC_47 NC_48 NC_49 NC_50 NC_51 NC_52 NC_53 Net-_U6-Pad17_ Net-_U6-Pad18_ Net-_U6-Pad19_ NC_54 Net-_U6-Pad21_ Net-_U6-Pad22_ NC_55 NC_56 MAX238
.end
