.title KiCad schematic
U1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 GND GND GND GND VCC GND GND GND GND VCC VCC NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 VCC VCC Net-_R1-Pad2_ NC_13 NC_14 GND Net-_R2-Pad2_ Net-_R3-Pad2_ Net-_R4-Pad2_ Net-_R5-Pad2_ Net-_R6-Pad2_ Net-_R7-Pad2_ Net-_R8-Pad2_ Net-_R9-Pad2_ NC_15 NC_16 NC_17 Z80ACPU
C1 VCC GND 1μF
R1 VCC Net-_R1-Pad2_ 470
SW1 GND Net-_R1-Pad2_ SW_SPST
R2 Net-_D1-Pad2_ Net-_R2-Pad2_ 330
R3 Net-_D2-Pad2_ Net-_R3-Pad2_ 330
R4 Net-_D3-Pad2_ Net-_R4-Pad2_ 330
R5 Net-_D4-Pad2_ Net-_R5-Pad2_ 330
R6 Net-_D5-Pad2_ Net-_R6-Pad2_ 330
R7 Net-_D6-Pad2_ Net-_R7-Pad2_ 330
R8 Net-_D7-Pad2_ Net-_R8-Pad2_ 330
R9 Net-_D8-Pad2_ Net-_R9-Pad2_ 330
D1 GND Net-_D1-Pad2_ LED
D2 GND Net-_D2-Pad2_ LED
D3 GND Net-_D3-Pad2_ LED
D4 GND Net-_D4-Pad2_ LED
D5 GND Net-_D5-Pad2_ LED
D6 GND Net-_D6-Pad2_ LED
D8 GND Net-_D8-Pad2_ LED
D7 GND Net-_D7-Pad2_ LED
.end
