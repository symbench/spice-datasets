.title KiCad schematic
K1 CTRL RZ03-1A4-D005
R4 NC_01 NC_02 R
R1 NC_03 NC_04 R
SW1 GND RST SW_PUSH_SMALL_H
IC1 RST NC_05 NC_06 NC_07 MOSI CTRL SCK NC_08 ATTINY85-S
P1 CTRL +5V SCK MOSI RST GND CONN_02X03
R2 NC_09 GND R
R3 NC_10 GND R
.end
