.title KiCad schematic
U1 NC_01 Net-_U1-Pad2_ NC_02 NC_03 NC_04 2SK2145-BL
U6 Net-_U6-Pad1_ Net-_U6-Pad1_ Net-_U6-Pad1_ NC_05 NC_06 NC_07 NC_08 Net-_U6-Pad10_ Net-_U6-Pad10_ Net-_U6-Pad10_ LT1995
U2 NC_09 Net-_U2-Pad2_ NC_10 NC_11 NC_12 2SK2145-BL
U7 Net-_U7-Pad1_ Net-_U7-Pad1_ Net-_U1-Pad2_ NC_13 NC_14 Net-_U2-Pad2_ DMMT3904
.end
