.title KiCad schematic
U3 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 DS1511Y+
J2 VCC VCC /D0 /A0 /D1 /A1 /D2 /A2 /D3 /A3 /D4 /A4 /D5 NC_26 /D6 NC_27 /D7 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 NC_43 NC_44 NC_45 NC_46 NC_47 NC_48 GND GND Expansion Bus
C5 GND VCC 0.1uF
U5 NC_49 NC_50 NC_51 NC_52 NC_53 /A4 /A3 /A2 /A1 /A0 /D0 /D1 /D2 GND /D3 /D4 /D5 /D6 /D7 NC_54 GND NC_55 GND NC_56 NC_57 NC_58 NC_59 VCC DS1501W
.end
