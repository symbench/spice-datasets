.title KiCad schematic
V1 vin 0 pulse(0 3.3 0 0 0 100m 200m)
V2 VDD 0 3.3
M1 vout vin VDD VDD MPMOS
M2 vout vin 0 0 MNMOS
.tran 1m 400m
.model mnmos nmos level=8 version=3.3.0
.model mpmos pmos level=8 version=3.3.0
.control
run
plot v(vin)+5 v(vout)
.endc
.end
