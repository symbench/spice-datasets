.title KiCad schematic
X1 Net-_C3-Pad1_ GND Net-_C4-Pad1_ GND 16MHz 18pF
C2 +12V GND 10uF 25V
C5 Net-_C5-Pad1_ GND 10uF 25V
C3 Net-_C3-Pad1_ GND 22pF
C4 Net-_C4-Pad1_ GND 22pF
D1 /VIN GND 14V
F1 +12V Net-_D2-Pad1_ 1.1A 25V
J1 /VIN GND INPUT
D2 Net-_D2-Pad1_ /VIN 20V 1A
C7 +5V GND 100nF
C8 +5V GND 100nF
C9 +5V GND 100nF
J3 /MISO2 +5V /SCK2 /MOSI2 /~RESET2 GND ISP-2560
U1 GND Net-_C5-Pad1_ +12V NCP1117-5V
C1 /~RESET2 /FTDI_RESET 100nF
J2 /FTDI_RESET /FTDI_TXOUT /FTDI_RXIN +5V NC_01 GND FTDI
D3 +5V Net-_C5-Pad1_ 20V 1A
LED1 GND NC_02 AMBER
C6 +5V GND 100nF
C10 +5V GND 100nF
U2 /FTDI_RXIN /FTDI_TXOUT +5V GND /SCK2 /MOSI2 /MISO2 NC_03 /~RESET2 +5V GND Net-_C3-Pad1_ Net-_C4-Pad1_ +5V GND +5V GND +5V GND +5V ATMEGA2560
S1 GND /~RESET2 RESET
.end
