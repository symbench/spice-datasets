.title KiCad schematic
XA1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 S0 S1 S2 S3 S4 S5 S6 NC_13 NC_14 NC_15 NC_16 NC_17 GND NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 +5V Arduino_Uno_Shield
SW6 GND S5 +5V SW_SPDT
SW5 GND S4 +5V SW_SPDT
SW4 GND S3 +5V SW_SPDT
SW3 GND S2 +5V SW_SPDT
SW2 GND S1 +5V SW_SPDT
SW1 GND S0 +5V SW_SPDT
SW7 GND S6 +5V SW_SPDT
.end
