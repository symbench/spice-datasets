.title KiCad schematic
J1 Net-_J1-Pad1_ Net-_J1-Pad2_ C
J2 Net-_J1-Pad1_ Net-_J1-Pad2_ C
J3 Net-_J1-Pad1_ Net-_J1-Pad2_ C
.end
