.title KiCad schematic
D1 +5V Net-_D1-Pad2_ LED
D2 +12V Net-_D2-Pad2_ LED
D3 Net-_D3-Pad1_ -12V LED
R1 Net-_D1-Pad2_ GND 270
R2 Net-_D2-Pad2_ GND 1k
R3 Net-_D3-Pad1_ GND 1k
J2 -12V -12V GND GND GND GND GND GND +12V +12V +5V +5V CV CV GATE GATE Conn_02x08_Row_Letter_Last
J10 -12V -12V GND GND GND GND GND GND +12V +12V +5V +5V CV CV GATE GATE Conn_02x08_Row_Letter_Last
J11 -12V -12V GND GND GND GND GND GND +12V +12V +5V +5V CV CV GATE GATE Conn_02x08_Row_Letter_Last
J12 -12V -12V GND GND GND GND GND GND +12V +12V +5V +5V CV CV GATE GATE Conn_02x08_Row_Letter_Last
J3 -12V -12V GND GND GND GND GND GND +12V +12V +5V +5V CV CV GATE GATE Conn_02x08_Row_Letter_Last
J5 -12V -12V GND GND GND GND GND GND +12V +12V +5V +5V CV CV GATE GATE Conn_02x08_Row_Letter_Last
J7 -12V -12V GND GND GND GND GND GND +12V +12V +5V +5V CV CV GATE GATE Conn_02x08_Row_Letter_Last
J9 -12V -12V GND GND GND GND GND GND +12V +12V +5V +5V CV CV GATE GATE Conn_02x08_Row_Letter_Last
J8 -12V -12V GND GND GND GND GND GND +12V +12V +5V +5V CV CV GATE GATE Conn_02x08_Row_Letter_Last
J13 -12V -12V GND GND GND GND GND GND +12V +12V +5V +5V CV CV GATE GATE Conn_02x08_Row_Letter_Last
J6 -12V -12V GND GND GND GND GND GND +12V +12V +5V +5V CV CV GATE GATE Conn_02x08_Row_Letter_Last
J4 -12V -12V GND GND GND GND GND GND +12V +12V +5V +5V CV CV GATE GATE Conn_02x08_Row_Letter_Last
J1 -12V GND +12V +5V CV GATE Screw_Terminal_01x06
.end
