.title KiCad schematic
U201 /JTAG_TCK NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 /JTAG_TDO /JTAG_TDI ~RESET NC_07 NC_08 NC_09 /JTAG_TMS COM NC_10 NC_11 NC_12 ONOFF NC_13 NC_14 NC_15 NC_16 Net-_J1102-Pad2_ Net-_C1104-Pad1_ Net-_C1101-Pad1_ Net-_C1102-Pad1_ NC_17 NC_18 Net-_C1103-Pad1_ MCIMX6Y2DVM
Y1101 Net-_C1101-Pad1_ COM Net-_C1102-Pad1_ COM 24MHz
C1102 Net-_C1102-Pad1_ COM 6p
C1101 Net-_C1101-Pad1_ COM 6p
Y1102 Net-_C1103-Pad1_ Net-_C1104-Pad1_ 32.768kHz
C1104 Net-_C1104-Pad1_ COM 19p
C1103 Net-_C1103-Pad1_ COM 19p
J1102 PP_SNVS_IN Net-_J1102-Pad2_ FORCE SERIAL
J1101 PP_GPIO /JTAG_TMS COM /JTAG_TCK COM /JTAG_TDO NC_19 /JTAG_TDI COM ~RESET JTAG
S1101 NC_20 COM NC_21 ONOFF TACTILE-4
S1102 NC_22 COM NC_23 ~RESET TACTILE-4
U1102 /JTAG_TDI COM /JTAG_TDO /JTAG_TMS PP_GPIO /JTAG_TCK NUP4114
U1101 ONOFF COM NC_24 ~RESET PP_SNVS_IN NC_25 NUP4114
.end
