.title KiCad schematic
R1 Net-_R1-Pad1_ Net-_C1-Pad1_ 1k
C1 Net-_C1-Pad1_ 0 10u
V1 Net-_R1-Pad1_ 0 pulse(0 5 10m 1u 1u 1m 2m)
.end
