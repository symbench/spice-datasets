.title KiCad schematic
N2 20190606
N1 OHWLOGO
.end
