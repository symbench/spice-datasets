.title KiCad schematic
U6 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 THS4032ID
U8 NC_09 NC_10 AVDD NC_11 NC_12 GND NC_13 NC_14 THS4551IDGKT
U7 NC_15 NC_16 AVDD NC_17 NC_18 GND NC_19 NC_20 THS4551IDGKT
J16 NC_21 GND NC_22 NC_23 NC_24 NC_25 GND MDD01
.end
