.title KiCad schematic
U1 NC_01 NC_02 GND +5V GND +5V NC_03 NC_04 NC_05 NC_06 Net-_R1-Pad2_ NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 GND NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 ATmega328-AU
J1 GND +5V Conn_01x02_Female
R1 Net-_D1-Pad2_ Net-_R1-Pad2_ 361
D1 GND Net-_D1-Pad2_ LED
R3 +5V Net-_R3-Pad2_ 1k
R2 Net-_D2-Pad1_ GND 360
D2 Net-_D2-Pad1_ Net-_D2-Pad2_ LED
SW1 GND Net-_SW1-Pad2_ Pulsador
J2 GND +5V Conn_01x02_Female
U2 Net-_R3-Pad2_ Net-_D2-Pad2_ Net-_SW1-Pad2_ NC_27 NC_28 NC_29 +5V GND NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 GND NC_43 NC_44 NC_45 NC_46 NC_47 NC_48 ATmega328-PU
.end
