.title KiCad schematic
U1 GND VOUT FB EN SW +BATT GND FAN4860
P1 +BATT SW EN FB VOUT GND CONN_01X06
.end
