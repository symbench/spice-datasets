.title KiCad schematic
U1 /A15 /A14 /A13 /A12 /A11 /A10 /A9 /A8 NC_01 NC_02 /~WE +3V3 NC_03 +3V3 GND /A18 /A17 /A7 /A6 /A5 /A4 /A3 /A2 /A1 /A0 GND GND /~OE /D0 NC_04 /D1 NC_05 /D2 NC_06 /D3 NC_07 +3V3 /D4 NC_08 /D5 NC_09 /D6 NC_10 /D7 /A19 GND GND /A16 CY62157
C1 GND +3V3 0.1uF
J1 +3V3 GND /D0 /D1 /D2 /D3 /D4 /D5 /D6 /D7 /~OE /~WE /A19 /A18 /A17 /A16 Conn_01x16_Male
J2 GND NC_11 /A0 /A1 /A2 /A3 /A4 /A5 /A6 /A7 /A8 /A9 /A10 /A11 /A12 /A13 /A14 /A15 Conn_01x18_Male
.end
