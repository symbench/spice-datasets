.title KiCad schematic
BT1 Net-_BT1-Pad1_ Net-_BT1-Pad2_ 9V
R1 Net-_D1-Pad1_ Net-_C1-Pad1_ 470R
R2 Net-_BT1-Pad1_ Net-_C1-Pad2_ 47K
R3 Net-_BT1-Pad1_ Net-_C2-Pad2_ 47K
R4 Net-_D2-Pad1_ Net-_C2-Pad1_ 470R
D1 Net-_D1-Pad1_ Net-_BT1-Pad1_ LED
D2 Net-_D2-Pad1_ Net-_BT1-Pad1_ LED
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 47uF
C2 Net-_C2-Pad1_ Net-_C2-Pad2_ 47uF
U1 Net-_BT1-Pad2_ Net-_C1-Pad2_ Net-_C1-Pad1_ Net-_BT1-Pad2_ Net-_C2-Pad2_ Net-_C2-Pad1_ BC846BDW1T1G
.end
