.title KiCad schematic
U1 Net-_J2-Pad4_ Net-_J2-Pad2_ X Net-_J2-Pad1_ Net-_J2-Pad3_ I E VSS C B A Net-_J2-Pad5_ Net-_J2-Pad8_ Net-_J2-Pad7_ Net-_J2-Pad6_ VDD 4051
U2 Net-_J2-Pad4_ Net-_J2-Pad2_ X Net-_J2-Pad1_ Net-_J2-Pad3_ I E VSS C B A Net-_J2-Pad5_ Net-_J2-Pad8_ Net-_J2-Pad7_ Net-_J2-Pad6_ VDD 4051
J2 Net-_J2-Pad1_ Net-_J2-Pad2_ Net-_J2-Pad3_ Net-_J2-Pad4_ Net-_J2-Pad5_ Net-_J2-Pad6_ Net-_J2-Pad7_ Net-_J2-Pad8_ Conn_01x08
J1 VDD X I E A B C VSS Conn_01x08
C1 VDD VSS C_Small
R1 I VSS 10K
.end
