.title KiCad schematic
J1 NC_01 NC_02 /FCR2_1 /FCR2_2 /FCU1_1 /FCU1_2 /FDP1_1 /FDP1_2 /FDS1_1 /FDS1_2 /FDP3_1 /FDP3_2 /PT_1 /PT_2 /APB_1 /APB_2 /FPB_1 /FPB_2 /Lum_1 /Lum_2 /fDI_1 /fDI_2 /SUP_1 /SUP_2 /ECU_1 /ECU_2 /ECR_2 /ECR_3 /EDC1_1 /EDC1_2 /BI_1 /BI_2 /TRI_1 /TRI_2 NC_03 /OmneticsRef Conn_02x18_Odd_Even
J2 /FDP2_1 /FDP2_2 /FCR2_1 /FCR2_2 /FCU1_1 /FCU1_2 /FCU2_1 /FCU2_2 /FCR1_1 /FCR1_2 /FDP1_1 /FDP1_2 /FDS1_1 /FDS1_2 /FDS2_1 /FDS2_2 /FDP3_1 /FDP3_2 /PT_1 /PT_2 /APB_1 /APB_2 /FPB_1 /FPB_2 /Lum_1 /Lum_2 /fDI_1 /fDI_2 NC_04 NC_05 /SUP_1 /SUP_2 /ECU_1 /ECU_2 NC_06 NC_07 /ECR_2 /ECR_3 /EDC1_1 /EDC1_2 /EDC2_1 /EDC2_2 /BI_1 /BI_2 /TRI_1 /TRI_2 /SamtecRef1 /SamtecRef2 /SamtecRef3 /SamtecRef4 Conn_02x25_Odd_Even
U1 /OmneticsRef /SamtecRef1 /SamtecRef2 /SamtecRef3 /SamtecRef4 SamtecReferences
J3 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 NC_43 NC_44 NC_45 NC_46 NC_47 NC_48 NC_49 NC_50 NC_51 NC_52 NC_53 /SamtecRef1 /SamtecRef2 /SamtecRef3 /SamtecRef4 Conn_02x25_Odd_Even
J4 NC_54 NC_55 /FDP2_1 /FDP2_2 /FCR2_1 /FCR2_2 /FCU1_1 /FCU1_2 /FCU2_1 /FCU2_2 /FCR1_1 /FCR1_2 /FDP1_1 /FDP1_2 /FDS1_1 /FDS1_2 /FDS2_1 /FDS2_2 /FDP3_1 /FDP3_2 /APB_1 /APB_2 /FPB_1 /FPB_2 /Lum_1 /Lum_2 /ECU_1 /ECU_2 /ECR_2 /ECR_3 /EDC1_1 /EDC1_2 /EDC2_1 /EDC2_2 NC_56 /OmneticsRef Conn_02x18_Odd_Even
U2 /OmneticsRef /SamtecRef1 /SamtecRef2 /SamtecRef3 /SamtecRef4 SamtecReferences
.end
