.title KiCad schematic
U1 GND Net-_C2-Pad2_ Measure1 Measure3.2 Net-_C1-Pad2_ Net-_C2-Pad2_ Net-_R1-Pad1_ VCC LM555N
C1 GND Net-_C1-Pad2_ 10n
R2 Net-_R1-Pad1_ Net-_C2-Pad2_ 12k
R1 Net-_R1-Pad1_ Measure3.2 2.2k
SW1 NC_01 VCC Net-_1N400X1-Pad2_ SWITCH_INV
1N400X1 VCC Net-_1N400X1-Pad2_ D
C7 VCC GND 220u
C8 /12V GND 47u
C9 Measure3.2 GND 47u
R5 Net-_D5-Pad2_ Measure3.2 270
D5 GND Net-_D5-Pad2_ LED
2N2222 Net-_2N2222-Pad1_ Net-_2N2222-Pad2_ GND Q_NPN_BCE
R4 VCC Net-_2N2222-Pad2_ 1.8k
2N2222_1 Net-_2N2222-Pad2_ VCC Measure2 Q_NPN_BCE
2N2907 Net-_2N2222-Pad2_ GND Measure2 Q_PNP_BCE
C3 Measure2 Net-_1N400X2-Pad2_ 47u
1N400X2 GND Net-_1N400X2-Pad2_ D
1N400X3 Net-_1N400X2-Pad2_ Net-_-12V1-PadVI_ D
C4 GND Net-_-12V1-PadVI_ 47u
C5 GND Net-_-12V1-PadVO_ 47u
R3 Net-_2N2222-Pad1_ Measure1 3.3k
C2 GND Net-_C2-Pad2_ 47n
-12V1 GND Net-_-12V1-PadVI_ Net-_-12V1-PadVO_ LM2990
-5V1 GND Net-_-12V1-PadVO_ /-5V LM2990
C6 GND /-5V 47u
+12V1 GND VCC /12V LM2940
+5V1 GND /12V Measure3.2 LM2940
.end
