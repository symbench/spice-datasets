.title KiCad schematic
IC1 Net-_IC1-Pad1_ Prog Net-_IC1-Pad3_ GND NEO Net-_IC1-Pad6_ Net-_IC1-Pad7_ VCC ATTINY85-20PU
R1 VCC Prog 22K
JACK1 GND NC_01 Net-_C1-Pad2_ NC_02 NC_03 NC_04 JACK_TRS_6PINS
JACK2 GND Net-_JACK2-Pad2_ NC_05 NC_06 NC_07 NC_08 JACK_TRS_6PINS
C1 Prog Net-_C1-Pad2_ 100nF
C2 GND VCC 100nF
R2 Prog GND 22K
R3 Prog Net-_PUSH1-Pad1_ 22K
PUSH1 Net-_PUSH1-Pad1_ GND SW_Push
SW1 +BATT VCC SW_SPST
R4 Net-_POT1-Pad2_ Net-_IC1-Pad7_ 22K
POT1 GND Net-_POT1-Pad2_ Net-_POT1-Pad3_ POT
R5 Net-_POT1-Pad3_ VCC 4K7
R6 Net-_IC1-Pad6_ Net-_D1-Pad2_ 1K
D1 GND Net-_D1-Pad2_ LED
TRIM1 Net-_C3-Pad2_ Net-_JACK2-Pad2_ GND POT
R7 Net-_C3-Pad2_ Net-_IC1-Pad6_ 330
C3 GND Net-_C3-Pad2_ 100nF
J6 Net-_IC1-Pad6_ PB1
J5 NEO PB0
J7 Net-_IC1-Pad7_ PB2
J2 Prog PB3
J3 Net-_IC1-Pad3_ PB4
J1 Net-_IC1-Pad1_ PB5
J4 GND GND
J8 VCC VCC
J9 Net-_C1-Pad2_ Prog
J10 Net-_C3-Pad2_ S-Out
J11 Net-_D1-Pad2_ LED
NEO2 VCC NC_09 GND Net-_NEO1-Pad2_ SK6813b
NEO1 VCC Net-_NEO1-Pad2_ GND NEO SK6813b
.end
