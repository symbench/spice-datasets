.title KiCad schematic
U1 Net-_R1-Pad2_ NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 /3.3V GND NC_07 NC_08 NC_09 NC_10 NC_11 /RXD NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 ESP-12E
R2 NC_19 /RXD 1K
SW1 Net-_R1-Pad2_ GND SW_Push
R1 /3.3V Net-_R1-Pad2_ 10k
U2 GND MIC5524
C2 /Voltage Regulation/3.3V GND 10uF
C1 /Voltage Regulation/VBUS GND 10uF
R3 /Voltage Regulation/VBUS /Voltage Regulation/EN 10k
P1 NC_20 NC_21 NC_22 NC_23 GND NC_24 USB_OTG
C3 NC_25 GND 5uF
P2 NC_26 NC_27 NC_28 /Connectors/GPIO14/SCK /Connectors/GPIO12/MISO /Connectors/GPIO13/MOSI NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 CONN_01X12
P3 NC_35 NC_36 NC_37 /Connectors/GPIO12/MISO /Connectors/GPIO13/MOSI /Connectors/GPIO14/SCK NC_38 NC_39 NC_40 NC_41 NC_42 NC_43 GND NC_44 NC_45 NC_46 CONN_01X16
.end
