.title KiCad schematic
R2 RPI_19 3.3V 10k
Q1 D7 3.3V RPI_19 BS170
R1 D7 5V 10k
R4 RPI_18 3.3V 10k
Q2 D6 3.3V RPI_18 BS170
R3 D6 5V 10k
R6 RPI_17 3.3V 10k
Q3 D5 3.3V RPI_17 BS170
R5 D5 5V 10k
R8 RPI_16 3.3V 10k
Q4 D4 3.3V RPI_16 BS170
R7 D4 5V 10k
R10 RPI_15 3.3V 10k
Q5 D3 3.3V RPI_15 BS170
R9 D3 5V 10k
R12 RPI_14 3.3V 10k
Q6 D2 3.3V RPI_14 BS170
R11 D2 5V 10k
R14 RPI_13 3.3V 10k
Q7 D1 3.3V RPI_13 BS170
R13 D1 5V 10k
R16 RPI_12 3.3V 10k
Q8 D0 3.3V RPI_12 BS170
R15 D0 5V 10k
R18 RPI_10 3.3V 10k
Q9 RPI_SEL 3.3V RPI_10 BS170
R17 RPI_SEL 5V 10k
.end
