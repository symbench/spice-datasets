.title KiCad schematic
U3 /RO /DE /DE /DI GND /A /B +3V3 MAX3485
U2 Net-_R2-Pad2_ NC_01 Net-_R1-Pad2_ NC_02 NC_03 NC_04 Net-_R5-Pad2_ +3V3 GND /DE NC_05 /FLASH /DI /RO /RX /TX ESP-12E
R2 +3V3 Net-_R2-Pad2_ 10k
R1 +3V3 Net-_R1-Pad2_ 10k
U1 /AC_L /AC_N GND +3V3 HLK-PM03
J1 /AC_N /L 220AC
R4 +3V3 /FLASH 10k
C3 +3V3 GND 470uF
C1 +3V3 GND 0.1uF
C2 +3V3 GND 0.01uF
R3 /DE GND 5.7k
F1 /AC_L /L 250mA
RV1 /AC_L /AC_N S14K385
J3 /A /B RS485
C4 GND +3V3 0.1uF
J2 /TX /RX GND GND /FLASH +3V3 Conn_01x06_Male
SW1 GND Net-_R2-Pad2_ Reset
R5 Net-_D1-Pad2_ Net-_R5-Pad2_ 680
D1 GND Net-_D1-Pad2_ LED
R7 /B /A 120
R6 GND /B 560
R8 /A +3V3 560
R9 +3V3 /RO 10k
.end
