.title KiCad schematic
P8 /BAT_INT GND CONN_BAT_INT
P9 GND /SCK0/FRAME_STOP /EP_TXD /EP_RXD CONN_EP_UART
P1 GND /UART_VCC /UART_TX /UART_RX /HOST_INT CONN_UART
P2 /SRV_CAM /SRV_VOUT GND CONN_SRV_CAM
P3 /SRV_LOCK /SRV_VOUT GND CONN_SRV_LOCK
P4 /SRV_BRAKE /SRV_VOUT GND CONN_SRV_BRAKE
P5 /SRV_FOOT /SRV_VOUT GND CONN_SRV_FOOT
P7 /FAN_PWM /FAN_TACHO /FAN_VOUT GND CONN_FAN
P15 /STEP_B1 /STEP_B2 /STEP_A2 /STEP_A1 CONN_STEP
P16 /EP_VCC /EP_VCC GND GND CONN_EP_VCC
P14 VCC VCC GND GND CONN_VCC
P12 /BUTTON GND CONN_BTN
P13 /LED_VOUT GND /LED_CLK /LED_DAT CONN_LED
P17 VCC /IR_TX /IR_RX GND CONN_IR
R1 /UART_VCC /UART_TX 100K
P20 /EP_RXD /UART_TX /EP_TXD /UART_RX /SRV_CAM /SRV_FOOT /SRV_BRAKE /SRV_LOCK /A2 /SRV_VOUT /MOSI0/STEP_STOP1 /MISO0/STEP_STOP2 /SCK0/FRAME_STOP CONN1
P18 /CHG2_STAT/MISO1 /CHG2_CTL/MOSI1 /BAT2_CTL/SCK1 /FAN_VOUT /TMP_INT /FAN_PWM /HOST_INT /FAN_TACHO /~RESET0 /SCL0 /SDA0 /BUTTON /LED_DAT /LED_CLK /LED_VOUT CONN2
P21 /STEP_A1 /STEP_A2 /STEP_B2 /STEP_B1 /EP_VCC /EP_VCC CONN3
P22 NC_01 /SDA1 /SCL1 /~RESET1 /IR_TX /IR_RX /BAT_INT /SDA0 /SCL0 CONN4
P19 GND VCC CONN_VCC
P6 GND /MOSI0/STEP_STOP1 /MISO0/STEP_STOP2 CONN_STEP_STOP
P11 /~RESET1 /BAT2_CTL/SCK1 /CHG2_CTL/MOSI1 /CHG2_STAT/MISO1 CONN_SPI1
P10 /SCK0/FRAME_STOP /MISO0/STEP_STOP2 /MOSI0/STEP_STOP1 /~RESET0 CONN_SPI0
TP4 /A2 TEST_1P
P23 /SDA0 /SCL0 CONN_I2C0
P24 /SDA1 /SCL1 CONN_I2C1
P25 /SDA0 /SCL0 CONN_I2C2
P26 GND /TMP_INT /SCL1 /SDA1 VCC CONN_TMP
.end
