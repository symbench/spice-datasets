.title KiCad schematic
U1 DRIVE BAT SENSE TIMER Vin GND PROG Vin Vin GND NC_01 GND NC_02 Vin ~CHRG GND GND LTC4060
U2 DRIVE SENSE BAT MJD210
R2 Vin Net-_D1-Pad2_ 330
D1 ~CHRG Net-_D1-Pad2_ LED
R3 PROG GND 698
C1 TIMER GND 1.5n
U4 Vin NC_03 NC_04 NC_05 GND 609-4613-6-ND
P1 GND BAT CONN_01X02
U3 BAT GND Net-_U3-Pad3_ Net-_U3-Pad3_ 36-1022-ND
.end
