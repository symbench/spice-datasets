.title KiCad schematic
BT1 /VCC GND Battery 3V
C1 GND Net-_C1-Pad2_ 22pF
C2 GND Net-_C2-Pad2_ 22pF
C3 /VCC GND 10uF
D1 Net-_D1-Pad1_ /SCK LED
R1 Net-_D1-Pad1_ GND 330Ohm
R2 /VCC /RESET 10kOhm
U1 /ADDS1 /ADDS2 /VCC GND /SDA /SCL GND /VCC 24LC1025
U4 /D3 /D4 GND /VCC GND /VCC Net-_C1-Pad2_ Net-_C2-Pad2_ /D5 /D6 /D7 /D8 NC_01 NC_02 /MOSI /MISO /SCK /VCC NC_03 /VCC GND NC_04 /ADDS1 /ADDS2 NC_05 NC_06 /SDA /SCL /RESET /RX /TX /D2 ATMEGA328P-AU
U3 Net-_U3-Pad1_ Net-_U3-Pad2_ /VCC GND /SDA /SCL NC_07 /VCC DS1337_v1
Y1 Net-_U3-Pad1_ Net-_U3-Pad2_ Crystal 32 MHz
Y2 Net-_C1-Pad2_ Net-_C2-Pad2_ Crystal 16 MHz
U2 /ADDS1 /ADDS2 /VCC GND /SDA /SCL GND /VCC 24LC1025
J2 /D2 /D3 /D4 /D5 /D6 /D7 /D8 GND /VCC Digital pins
J4 GND /VCC /SDA /SCL I2C
J3 /MISO /VCC /SCK /MOSI /RESET GND ICSP
J1 GND /VCC /RX /TX Serial
.end
