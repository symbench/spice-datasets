.title KiCad schematic
J4 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 Conn_02x03_Male_ICSP
.end
