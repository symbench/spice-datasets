.title KiCad schematic
UK12 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 /RTC-O /RTC-CLK /RTC-CS* ADB-INT* ADB-ST0 ADB-ST1 NC_09 NC_10 ADB-SCLK ADB-DIO NC_11 R-W* NC_12 PU E /D_31_ /D_30_ /D_29_ /D_28_ /D_27_ /D_26_ /D_25_ /D_24_ RESET* /A_12_ /A_11_ /A_10_ /A_9_ /RTC-1HZ VBLK* 65C22
UK11 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 VBLK* NC_28 NC_29 NC_30 R-W* NC_31 PU E /D_31_ /D_30_ /D_29_ /D_28_ /D_27_ /D_26_ /D_25_ /D_24_ RESET* /A_12_ /A_11_ /A_10_ /A_9_ NC_32 NC_33 65C22
UL11 NC_34 /ADB0 /ADB0 RESET* NC_35 NC_36 ADB-SCLK ADB-DIO ADB-INT* NC_37 NC_38 NC_39 NC_40 ADB-ST0 ADB-ST1 ADB
J9 Net-_J9-Pad~_ ADB_CONN
J10 /ADBF ADB_CONN
L1 NC_41 /ADB0 NC_42 NC_43 /GNDF-ADB /+5F-ADB /ADBF NC_44 LNET
BT1 Button
UK4 /RTC-1HZ NC_45 NC_46 NC_47 /RTC-CS* /RTC-O /RTC-CLK NC_48 RTC
.end
