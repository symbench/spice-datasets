.title KiCad schematic
J3 Net-_FB2-Pad2_ Net-_J2-Pad1_ Net-_J1-Pad2_ NC_01 GND 10118194-0001LF
C9 GND +5V 10uF
FB2 +5V Net-_FB2-Pad2_ 1A 50m
J2 Net-_J2-Pad1_ NC_02 61300211121
J1 NC_03 Net-_J1-Pad2_ 61300211121
U1 NC_04 NC_05 NC_06 NC_07 NC_08 AP3429A
.end
