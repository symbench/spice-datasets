.title KiCad schematic
J1 +5V NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 GND Conn_01x12
.end
