.title KiCad schematic
J1 GND NC_01 NC_02 NC_03 /15V_UnProtected GND /PIC32_RX /PIC32_~RX /PIC32_~TX /PIC32_TX DB9_Female_MountingHoles
U1 +9V GND +5V L7805
U?1 +5V /ESP32_RX_5V NC_04 GND /PIC32_RX /PIC32_~RX /PIC32_~TX /PIC32_TX SN75179BD
R1 Net-_D3-Pad2_ /ESP32_RX_5V 1K
D3 +3V3 Net-_D3-Pad2_ 1N4148
D6 Net-_D6-Pad1_ NC_05 LED
D5 Net-_D5-Pad1_ NC_06 LED
R3 Net-_D5-Pad1_ GND 220
R4 Net-_D6-Pad1_ GND 220
U3 Net-_C1-Pad1_ GND +9V L7809
C2 +9V GND 0.1uF 16V
C3 +5V GND 0.1uF 16V
C1 Net-_C1-Pad1_ GND 0.33uF 50v
J2 +3V3 +5V +9V GND NC_07 NC_08 Conn_01x06_Female
D1 Net-_C1-Pad1_ /15V_UnProtected B120-E3
D2 GND Net-_D2-Pad2_ LED
R2 +5V Net-_D2-Pad2_ 470
U2 Net-_U2-Pad1_ NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 Net-_U2-Pad1_ NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 NC_43 Net-_U2-Pad1_ ESP32-WROOM-32D
.end
