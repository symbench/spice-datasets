.title KiCad schematic
P3 /VOUT NC_01 GND CONN_01X01
C1 /V5 GND 1uF
C2 /BAT GND 22uF
R2 Net-_R1-Pad2_ GND 30.1K
C3 /VOUT GND 22uF
R1 /VOUT Net-_R1-Pad2_ 102K
P1 GND /BAT /V5 CONN_01X01
.end
