.title KiCad schematic
R3 Net-_C1-Pad1_ GND 150R
C1 Net-_C1-Pad1_ L_OUT 47uF
C2 Net-_C2-Pad1_ R_OUT 47uF
R4 GND Net-_C2-Pad1_ 150R
C3 Net-_C1-Pad1_ GND 33nF
C4 GND Net-_C2-Pad1_ 33nF
R5 L_IN_FIL Net-_C1-Pad1_ 270R
R6 R_IN_FIL Net-_C2-Pad1_ 270R
U2 Net-_R10-Pad2_ GND Net-_R7-Pad2_ L_IN_FIL +3V3 R_IN_FIL NC7WZ16
R1 L_OUT GND 1.8K
R2 GND R_OUT 1.8K
R9 L_IN_UNF Net-_R7-Pad2_ 100R
R10 R_IN_UNF Net-_R10-Pad2_ 100R
R7 GND Net-_R7-Pad2_ 470R
R8 GND Net-_R10-Pad2_ 470R
U1 VCC GND VCC Net-_C5-Pad1_ +3V3 MIC5219-3.3BM5
C5 Net-_C5-Pad1_ GND 470pF
C6 +3V3 GND 2.2uF
TP1 L_OUT L_OUT
TP3 R_OUT R_OUT
TP4 L_IN_FIL LIN_FIL
TP6 R_IN_FIL RIN_FIL
TP7 L_IN_UNF LIN_RAW
TP9 R_IN_UNF RIN_RAW
TP10 +3V3 3V3
TP11 GND GND
TP5 GND GND
TP2 GND GND
TP8 GND GND
TP12 VCC VIN
C7 +3V3 GND 100nF
.end
