.title KiCad schematic
U1 OUT2 OUT1 +BATT BAT_SENSE Net-_RN1-Pad2_ BAT_SENSE Net-_RN1-Pad3_ BAT_SENSE Net-_RN1-Pad5_ BAT_SENSE Net-_RN1-Pad4_ GND OUT3 OUT4 LM339
D1 GND REF 0
C1 +BATT GND 100nF
RN1 REF Net-_RN1-Pad2_ Net-_RN1-Pad3_ Net-_RN1-Pad4_ Net-_RN1-Pad5_ Net-_RN1-Pad4_ Net-_RN1-Pad3_ Net-_RN1-Pad2_ 1K
RN3 +BATT +BATT BAT_SENSE BAT_SENSE GND Net-_RN3-Pad6_ Net-_RN3-Pad6_ Net-_RN3-Pad6_ 10K
RN2 Net-_RN1-Pad5_ Net-_RN1-Pad5_ REF REF +BATT +BATT GND GND 10K
RN5 OUT1 OUT2 OUT3 OUT4 +BATT +BATT +BATT +BATT 10K
D2 GND Net-_D2-Pad2_ 1
D3 GND Net-_D3-Pad2_ 2
D4 GND Net-_D4-Pad2_ 3
D5 GND Net-_D5-Pad2_ 4
RN4 OUT1 OUT2 OUT3 OUT4 Net-_D5-Pad2_ Net-_D4-Pad2_ Net-_D3-Pad2_ Net-_D2-Pad2_ 1K
J2 OUT1 OUT2 OUT3 OUT4 Conn_01x04
J1 +BATT +BATT GND GND Conn_01x04
.end
