.title KiCad schematic
U1 /VCCA /VCCA Net-_J1-Pad2_ GND Net-_U1-Pad5_ /DAC2 /DAC2 +5V MC4558CPT
C1 GND +5V 0.1uF
U2 /DAC3 /DAC3 Net-_U2-Pad3_ GND Net-_U2-Pad5_ /DAC4 /DAC4 +5V MC4558CPT
C2 GND +5V 0.1uF
U3 +5V Net-_J1-Pad2_ Net-_U1-Pad5_ Net-_U2-Pad3_ Net-_U2-Pad5_ GND +5V NC_01 /SSEL NC_02 DAC084S085
R1 +5V /SSEL 10k
J1 GND Net-_J1-Pad2_ Conn_01x02_Female
U4 VCC GND VCC NC_03 +1V2 MIC94310
C4 +1V2 GND 10uF
C3 GND VCC 0.47uF
U5 VCC GND VCC NC_04 +2V5 MIC94310
C6 +2V5 GND 10uF
C5 GND VCC 0.47uF
.end
