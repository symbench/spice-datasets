.title KiCad schematic
U1 NC_01 Net-_R1-Pad2_ GND -12V NC_02 /AD0 +12V NC_03 OP07
R1 /SNS Net-_R1-Pad2_ R
U2 NC_04 /AD0 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 PIC18F452-IP
R2 Net-_R1-Pad2_ /AD0 R
J1 GND /SNS Screw_Terminal_01x02
.end
