.title KiCad schematic
U2 RST ADC CH_PD NC_01 UV_INT RTS CTS +3V3 GND GPIO15 BT_EN GPIO0 SDA SCL ESP_RXD ESP_TXD ESP-12
U1 GND +3V3 +VSW AZ1117-3.3
C1 VBUS GND 100nF
C2 +3V3 GND 10uF
C3 +3V3 GND 100nF
SW1 RST GND RST
SW2 GPIO0 GND GP0
J2 RTS BT_RXD BT_TXD +3V3 CTS GND BLUETOOTH
R5 +3V3 SDA 10K
R4 +3V3 SCL 10K
D1 +VSW VBUS D_Schottky
J1 VBUS NC_02 NC_03 NC_04 NC_05 NC_06 USB_OTG
U3 BT_EN BT_TXD ESP_RXD BT_EN ESP_TXD BT_RXD GND NC_07 GND Net-_R7-Pad2_ NC_08 GND Net-_R7-Pad2_ VCC 74125
R7 +3V3 Net-_R7-Pad2_ 10K
D2 +VSW +BATT D_Schottky
R1 +3V3 GPIO0 10K
R2 GND GPIO15 10K
R3 +3V3 BT_EN 10K
C5 +VSW GND 100nF
C4 +VSW GND 10uF
U4 GND UV_INT SDA Net-_R8-Pad1_ SCL +3V3 VEML6070
R6 +3V3 UV_INT 10K
R8 Net-_R8-Pad1_ GND 300K
C6 +3V3 GND 100nF
U5 VBUS GND +BATT GND TP4056_BREAKOUT
R9 +3V3 RST 10K
R10 +3V3 CH_PD 10K
J3 GND ADC EXT_WATER_SENSOR
RV1 ADC +3V3 +3V3 47K
C7 ADC GND 1nF
.end
