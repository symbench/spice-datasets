.title KiCad schematic
C19 +3V3 GND 10uF
SW2 GND /RST_BT BT_RST
RP12 +3V3 /RST_BT 10k
D2 /P2_7 Net-_D2-Pad2_ BT_TX_LED
RP11 Net-_D2-Pad2_ +3V3 1k
RP10 Net-_D1-Pad2_ +3V3 1k
D1 /P0_2 Net-_D1-Pad2_ BT_PLED
U7 NC_01 GND NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 /P0_2 GND +3V3 /P2_7 NC_11 RN4871-V/RM118
.end
