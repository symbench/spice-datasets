.title KiCad schematic
J1 GNDREF /VBAT+ 36V Battery
D10 Net-_C13-Pad1_ /VBAT+ 1N5061
U5 /12V_IR GNDREF GNDREF GNDREF Net-_C13-Pad1_ Net-_D11-Pad1_ LM2574HVM-12
C13 Net-_C13-Pad1_ GNDREF 100uF
L1 Net-_D11-Pad1_ /12V_IR 300uH
D11 Net-_D11-Pad1_ GNDREF 1N5828
C14 /12V_IR GNDREF 330uF
U6 /12V GNDREF /5V L7805
C15 /12V GNDREF CP1
C16 /5V GNDREF 0.1uF
U7 /12V Net-_C17-Pad2_ Net-_C17-Pad2_ Net-_C17-Pad2_ Net-_C17-Pad1_ Net-_D12-Pad1_ LM2574HVM-12
C17 Net-_C17-Pad1_ Net-_C17-Pad2_ 100uF
L2 Net-_D12-Pad1_ /12V 300uH
D12 Net-_D12-Pad1_ Net-_C17-Pad2_ 1N5828
C19 /12V Net-_C17-Pad2_ 330uF
U8 /3v3 Net-_C18-Pad2_ /5V LP2950-3.3_TO92
C18 /5V Net-_C18-Pad2_ 0.1uF
C20 /3v3 Net-_C18-Pad2_ 2.2uF
.end
