.title KiCad schematic
U1 VCC GND +5V GND BEC
C1 +5V GND 10u
J1 IO25=SPORT GND VCC /HEART_BEAT /PXX_OUT NC_01 NC_02 NC_03 Conn_XLite
C2 +3V3 GND 10u
C3 +3V3 GND 100u
U3 GND +3V3 +3V3 NC_04 NC_05 IO34=DIO0 IO35=MISO IO32=SCK IO33=HEART_BEAT_3V3 IO25=SPORT IO26=PXX_OUT_3V3 IO27=SCREEN_SCL IO14=SCREEN_SDA IO12=RGBLED GND IO13=RST NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 IO0=SW1 IO4=DIO5 IO16=DIO4 IO17=DIO3 IO5=DIO2 IO18=DIO1 IO19=MOSI NC_14 IO21=NSS RX0 TX0 IO22=TXEN IO23=RXEN GND GND ESP32-WROOM
SW1 GND IO0=SW1 SW_Push
J3 GND +3V3 IO27=SCREEN_SCL IO14=SCREEN_SDA Screen
U2 GND +3V3 +5V AMS1117-3.3
D1 /LED_RGB_5V NC_15 GND IO12=RGBLED WS2812B
R5 +5V /LED_RGB_5V 75
C4 /LED_RGB_5V GND 100n
U4 GND IO4=DIO5 IO16=DIO4 IO17=DIO3 IO5=DIO2 IO18=DIO1 IO34=DIO0 IO13=RST GND GND +5V IO32=SCK IO35=MISO IO19=MOSI IO21=NSS IO22=TXEN IO23=RXEN GND /ANT GND GND GND E19-XXXM30S
J2 GND TX0 RX0 Programming
AE1 /ANT GND Antenna_Dipole
Q1 +3V3 IO33=HEART_BEAT_3V3 /HEART_BEAT Q_NMOS_GSD
R1 VCC /HEART_BEAT 10k
R2 +3V3 IO33=HEART_BEAT_3V3 10k
Q2 +3V3 IO26=PXX_OUT_3V3 /PXX_OUT Q_NMOS_GSD
R3 VCC /PXX_OUT 10k
R4 +3V3 IO26=PXX_OUT_3V3 10k
.end
