.title KiCad schematic
U1 WORKING_1 NC_01 NC_02 REFERENCE COUNTER WORKING_6 SPEC
U2 WORKING_1 WORKING_6 SMM-102-02-S-S
U3 NC_03 NC_04 SMM-102-02-S-S
U4 COUNTER REFERENCE SMM-102-02-S-S
P1 REFERENCE COUNTER WORKING_6 WORKING_1 CONN_01X04
.end
