.title KiCad schematic
J1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 Conn_02x05_Top_Bottom
U1 GND +3V3 Net-_C5-Pad1_ LM1117-3.3
C3 +5V_BUS GND 100uF
C4 +5V_BUS GND 100uF
C1 +5V_BUS GND 100uF
C2 +5V_BUS GND 100uF
C7 +3V3 GND 100pF
C8 +3V3 GND 10uF
C9 +3V3 GND 10uF
C6 Net-_C5-Pad1_ GND 25V 10uF
C5 Net-_C5-Pad1_ GND 50V 100pF
.end
