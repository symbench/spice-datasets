.title KiCad schematic
K4 /PWM2 +5V GND CONN_3
K3 /D2 +5V GND CONN_3
K2 /PWM1 +5V GND CONN_3
K1 /D1 +5V GND CONN_3
R1 Net-_D1-Pad2_ GND 1k
D1 +5V Net-_D1-Pad2_ LED
P1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 +5V GND NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 /D1 NC_17 NC_18 /PWM1 Net-_P1-Pad23_ NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 /D2 /PWM2 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 CONN_20X2
.end
