.title KiCad schematic
P1 Net-_P1-Pad1_ NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 Net-_P1-Pad12_ NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 CONN_01X19
P2 Net-_P2-Pad1_ Net-_P2-Pad2_ NC_18 NC_19 NC_20 Net-_P2-Pad6_ NC_21 Net-_P2-Pad8_ NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 CONN_01X19
U1 Net-_P1-Pad12_ Net-_P1-Pad1_ Net-_P2-Pad2_ Net-_P2-Pad6_ Net-_P2-Pad8_ Net-_P2-Pad1_ PYB30
.end
