.title KiCad schematic
U3 GND +3V3 NC_01 NC_02 NC_03 Net-_R2-Pad1_ Net-_R3-Pad1_ NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 GND NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 GND GND ESP32-WROOM-32
D1 GND Net-_D1-Pad2_ LED
SW1 Net-_R1-Pad1_ +5V SW_Push
J1 +5V NC_33 NC_34 NC_35 GND NC_36 USB_B_Micro
C1 +5V GND C
U1 GND +3V3 +5V AMS1117-3.3
C2 +3V3 GND CP1
R1 Net-_R1-Pad1_ Net-_D1-Pad2_ 1000
J2 Net-_J2-PadR1_ Net-_J2-PadR1_ NC_37 NC_38 Net-_J2-PadS1_ Net-_J2-PadS1_ NC_39 NC_40 GND GND NC_41 NC_42 AudioJack3_Dual_Switch
U2 Net-_R3-Pad1_ Net-_R3-Pad2_ Net-_J2-PadS1_ GND Net-_J2-PadS1_ Net-_R2-Pad2_ Net-_R2-Pad1_ +3V3 LM358
R2 Net-_R2-Pad1_ Net-_R2-Pad2_ 10k
R3 Net-_R3-Pad1_ Net-_R3-Pad2_ 10k
R5 Net-_R3-Pad2_ GND 1k
R4 GND Net-_R2-Pad2_ 1k
.end
