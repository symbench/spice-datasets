.title KiCad schematic
U2 GND Net-_U2-Pad2_ Net-_U2-Pad3_ NC_01 NC_02 Net-_J5-Pad2_ Net-_J5-Pad3_ Net-_J4-Pad2_ Net-_J4-Pad3_ Net-_J3-Pad2_ Net-_J3-Pad3_ Net-_C75-Pad2_ +3V3 Net-_R9-Pad1_ NC_03 NC_04 +3V3 Net-_R5-Pad1_ +3V3 VBUS +3V3 Net-_D69-Pad1_ Net-_R13-Pad2_ Net-_R10-Pad2_ NC_05 +3V3 NC_06 Net-_C75-Pad2_ FE1.1s
D74 Net-_D69-Pad1_ Net-_D74-Pad2_ Green
D75 Net-_D74-Pad2_ Net-_D69-Pad1_ Green
D73 Net-_D69-Pad2_ Net-_D69-Pad1_ Green
D69 Net-_D69-Pad1_ Net-_D69-Pad2_ Green
R13 Net-_D74-Pad2_ Net-_R13-Pad2_ 330
R10 Net-_D69-Pad2_ Net-_R10-Pad2_ 330
D76 Net-_D76-Pad1_ Net-_D69-Pad1_ Red
R14 GND Net-_D76-Pad1_ 330
Y1 Net-_U2-Pad2_ Net-_U2-Pad3_ 12MHz
C3 GND VBUS 0.1uF
C74 GND VBUS 10uF
R5 Net-_R5-Pad1_ GND 100K
R9 Net-_R9-Pad1_ GND 2K7
C75 GND Net-_C75-Pad2_ 10uF
C76 GND Net-_C75-Pad2_ 0.1uF
C77 GND +3V3 0.1uF
C78 GND +3V3 10uF
R8 Net-_R5-Pad1_ VBUS 47K
J3 VBUS Net-_J3-Pad2_ Net-_J3-Pad3_ GND GND USB_A
J4 VBUS Net-_J4-Pad2_ Net-_J4-Pad3_ GND GND USB_A
J5 VBUS Net-_J5-Pad2_ Net-_J5-Pad3_ GND GND USB_A
.end
