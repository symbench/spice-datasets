.title KiCad schematic
R1 Net-_R1-Pad1_ 0 1k
R3 Net-_R3-Pad1_ Net-_R3-Pad2_ 833
R2 Net-_R2-Pad1_ Net-_R1-Pad1_ 5k
V1 Net-_R3-Pad2_ 0 sin(0 10 50 0)
V2 Net-_U1-Pad5_ 0 +15v
V3 Net-_U1-Pad4_ 0 -15v
U1 Net-_R3-Pad1_ Net-_R1-Pad1_ Net-_R2-Pad1_ Net-_U1-Pad4_ Net-_U1-Pad5_ OPAMP
.end
