.title KiCad schematic
C1201 GNDD +5V 100n
U1202 GNDD NC_01 /XA4 NC_02 /XA5 NC_03 /XA6 NC_04 NC_05 GNDD GNDD /XA3 NC_06 /XA2 NC_07 /XA1 NC_08 /XA0 GNDD +5V 74HC244
U1203 NC_09 /XD7 /XD6 /XD5 /XD4 /XD3 /XD2 /XD1 /XD0 GNDD NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 +5V 74HC245
U1201 /~XCD0 /~XIRQ0 /~IOCS0 /~XCD1 /~XIRQ1 /~IOCS1 /~XCD2 /~XIRQ2 /~IOCS2 /~XCD3 GNDD /~XIRQ3 /~IOCS3 /~XCD4 /~XIRQ4 /~IOCS4 NC_19 NC_20 +5V XIOCON_PDIP
J1201 +5V +5V /~XIRQ0 /~XIRQ1 /~XIRQ2 /~XIRQ3 /~XIRQ4 /XA0 /XA1 /XA2 /XA3 /XA4 /XA5 /XA6 /XD0 /XD1 /XD2 /XD3 /XD4 /XD5 /XD6 /XD7 NC_21 +5V +5V +5V +5V NC_22 NC_23 /~IOCS4 /~IOCS3 /~IOCS2 /~IOCS1 /~IOCS0 GNDD GNDD GNDD GNDD GNDD GNDD GNDD GNDD GNDD /~XCD4 /~XCD3 /~XCD2 /~XCD1 /~XCD0 +5V +5V Conn_02x25_Counter_Clockwise
C1204 +5V GNDD 100n
C1205 +5V GNDD 1u
C1202 +5V GNDD 100n
C1203 GNDD +5V 100n
RN1201 +5V /~XCD4 /~XCD3 /~XCD2 /~XCD1 /~XCD0 47k
.end
