.title KiCad schematic
J1 GND 5V Net-_J1-Pad3_ Net-_J1-Pad4_ L_EN R_EN L_PWM R_PWM CONN_02X04
U1 NC_01 L_IS RXD2 CHAN_A CHAN_B L_PWM R_PWM L_EN R_EN SCL2 SDA2 NC_02 NC_03 GND 5V NC_04 GND NC_05 NC_06 NC_07 SCK2 SCK1 NC_08 TXD2 TXD1 Net-_D1-Pad2_ NC_09 NC_10 MOSI2 MOSI1 ESP32-DEVKIT-V1
D1 Net-_D1-Pad1_ Net-_D1-Pad2_ LED
R1 Net-_J1-Pad3_ L_IS 10k
R2 RXD2 Net-_J1-Pad4_ 10k
C2 RXD2 NC_11 0.1µ
J2 GND Net-_J2-Pad2_ Net-_J2-Pad3_ 5V CONN_01X04
R3 CHAN_B Net-_J2-Pad3_ 10k
R4 CHAN_A Net-_J2-Pad2_ 10k
C1 L_IS GND 0.1µ
R5 5V Net-_J2-Pad3_ 10K
R6 5V Net-_J2-Pad2_ 10K
R7 Net-_D1-Pad1_ 5V R
C3 5V GND CP
CON1 5V GND CHAN_A MOSI1 NC_12 SCK1 L_EN R_EN L_PWM TXD1 UEXT-5V
CON2 5V GND CHAN_B MOSI2 RXD2 SCK2 SCL2 SDA2 R_PWM TXD2 UEXT-5V
.end
