.title KiCad schematic
J1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 Conn_01x10_Male
U2 +3V3 Net-_R1-Pad1_ Net-_R2-Pad1_ Net-_R3-Pad1_ Net-_R4-Pad1_ Net-_R5-Pad1_ Net-_R6-Pad1_ GND_C GND_I Net-_R12-Pad2_ Net-_R11-Pad2_ Net-_R10-Pad2_ Net-_R9-Pad2_ Net-_R8-Pad2_ Net-_R7-Pad2_ 3V3_I SI8661AB-B-IS1
U1 NC_11 GND_C CS2_W CS1_W NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 CLK_W MISO_W MOSI_W CS0_W NC_19 WeMos_mini
J2 +3V3 GND_C CS2_E CS0_E CLK_E MISO_E MOSI_E CS1_E GND_I 3V3_I CONN_01X10
C1 3V3_I GND_I 100nF
C2 +3V3 GND_C 100nF
R1 Net-_R1-Pad1_ CLK_W 50R
R2 Net-_R2-Pad1_ MOSI_W 50R
R3 Net-_R3-Pad1_ CS0_W 50R
R4 Net-_R4-Pad1_ CS1_W 50R
R5 Net-_R5-Pad1_ CS2_W 50R
R6 Net-_R6-Pad1_ MISO_W 50R
R7 CLK_E Net-_R7-Pad2_ 50R
R8 MOSI_E Net-_R8-Pad2_ 50R
R9 CS0_E Net-_R9-Pad2_ 50R
R10 CS1_E Net-_R10-Pad2_ 50R
R11 CS2_E Net-_R11-Pad2_ 50R
R12 MISO_E Net-_R12-Pad2_ 50R
MS1 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 NC_43 NC_44 NC_45 NC_46 NC_47 ADAFRUIT_FEATHERWING_FitHome
.end
