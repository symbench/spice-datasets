.title KiCad schematic
H1 MountingHole
H2 MountingHole
.end
