.title KiCad schematic
U3 Net-_R3-Pad2_ GND /+12V_IN_ADC_OUT /+12V_IN_ADC_OUT +3V3 LM321
U1 NC_01 GND NC_02 NC_03 +3V3 LM321
C2 +3V3 GND 0.1uf
U2 Net-_R1-Pad2_ GND /+5V_IN_ADC_OUT /+5V_IN_ADC_OUT +3V3 LM321
C1 +3V3 GND 0.1uf
U5 Net-_R7-Pad2_ GND /+12V_BUS_ADC_OUT /+12V_BUS_ADC_OUT +3V3 LM321
C4 +3V3 GND 0.1uf
U4 Net-_R5-Pad2_ GND /+5V_BUS_ADC_OUT /+5V_BUS_ADC_OUT +3V3 LM321
C3 +3V3 GND 0.1uf
R3 NC_04 Net-_R3-Pad2_ 10K
R4 Net-_R3-Pad2_ GND 3.3K
R7 NC_05 Net-_R7-Pad2_ 10K
R8 Net-_R7-Pad2_ GND 3.3K
R5 NC_06 Net-_R5-Pad2_ 3K
R6 Net-_R5-Pad2_ GND 4.7K
R1 NC_07 Net-_R1-Pad2_ 3K
R2 Net-_R1-Pad2_ GND 4.7K
.end
