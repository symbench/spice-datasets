.title KiCad schematic
U4 +3V3 CC_SCL0 +3V3 CC_SDA0 Net-_R16-Pad2_ Net-_R16-Pad2_ Net-_R14-Pad2_ Net-_R14-Pad2_ NC_01 NC_02 NC_03 NC_04 NC_05 GND GND GND GND GND GND GND Net-_C29-Pad1_ +3V3 +3V3 Net-_C30-Pad1_ LSM9DS1
C30 Net-_C30-Pad1_ GND 0.1uF
C29 Net-_C29-Pad1_ GND 0.01uF
R14 +3V3 Net-_R14-Pad2_ 10k
R16 +3V3 Net-_R16-Pad2_ 10k
C34 +3V3 GND 10uF
C33 +3V3 GND 0.1uF
C31 +3V3 GND 0.1uF
C36 +3V3 GND 0.1uF
C35 +3V3 GND 4.7uF
R19 Net-_R19-Pad1_ +3V3 100K
R11 +3V3 CC_SCL0 4.7k
R12 +3V3 CC_SDA0 4.7k
U6 GND Net-_R19-Pad1_ CC_SDA0 CC_SCL0 GND +3V3 GND +3V3 BMP280
.end
