.title KiCad schematic
U101 NC_01 NC_02 NC_03 NC_04 3V LP2980IM5-3.0/NOPB
U201 NC_05 Net-_PD201-Pad2_ VGND 3V VGND Net-_PD301-Pad2_ NC_06 NC_07 Net-_PD401-Pad2_ VGND NC_08 VGND Net-_PD501-Pad2_ NC_09 MCP6404
PD201 VGND Net-_PD201-Pad2_ VBPW34SR
PD301 VGND Net-_PD301-Pad2_ VBPW34SR
PD401 VGND Net-_PD401-Pad2_ VBPW34SR
PD501 VGND Net-_PD501-Pad2_ VBPW34SR
.end
