.title KiCad schematic
U3 NC_01 GND Net-_RV2-Pad2_ GND /386out +12V NC_02 NC_03 LM386
C3 Net-_C3-Pad1_ Net-_C3-Pad2_ 10uF
R3 Net-_R3-Pad1_ Net-_C3-Pad1_ 1k
R4 /741out Net-_R3-Pad1_ 220k
R7 Net-_C6-Pad2_ GND 10
RV2 AC Net-_RV2-Pad2_ GND 100k
D2 GND Net-_C2-Pad1_ 1N4148
D1 Net-_C2-Pad1_ Net-_C4-Pad1_ 1N4148
C6 /386out Net-_C6-Pad2_ 47nF
C2 Net-_C2-Pad1_ /741out 0.1uF
R1 +180V Net-_R1-Pad2_ 470k
C5 /386out Net-_C5-Pad2_ 1000uF
LS1 Net-_C5-Pad2_ GND 8
T1 Net-_C4-Pad1_ GND NC_04 GND Net-_R5-Pad2_ NC_05 Net-_R1-Pad2_ NC_06 +180V EM80
C4 Net-_C4-Pad1_ GND 0.1uF
R5 Net-_R5-Pad1_ Net-_R5-Pad2_ 3W 10
R6 +12V Net-_R5-Pad1_ 3W 10
RV1 AC Net-_C3-Pad2_ GND 100k
C1 +12V GND 0.1uF
U1 +12V NC_07 GND +180V GND NCH6100HV
U2 NC_08 Net-_R3-Pad1_ GND GND NC_09 /741out +12V NC_10 LM741
R2 AC GND 1k
J1 AC AC GND AC AC AudioJack3_SwitchTR
J2 +12V GND GND Barrel_Jack_Switch
C7 +180V GND 1uF
.end
