.title KiCad schematic
U6 Net-_U3-Pad12_ NC_01 Net-_U3-Pad2_ Net-_U3-Pad13_ NC_02 Net-_Q1-Pad2_ Net-_U6-PadJ1.8_ NC_03 Net-_U3-Pad3_ Net-_U6-PadJ5.2_ NC_04 Net-_U6-PadJ5.4_ NC_05 Net-_U6-PadJ5.3_ NC_06 Net-_U6-PadJ5.1_ NC_07 NC_08 NC_09 NC_10 NC_11 Net-_U6-PadJ113_ Net-_Q2-Pad1_ Net-_Q3-Pad1_ NC_12 Net-_U3-Pad9_ Net-_R5-Pad1_ NC_13 NC_14 NC_15 NC_16 Net-_U6-PadJ512_ Net-_U6-PadJ513_ NC_17 NC_18 Net-_U6-PadJ516_ Net-_U6-PadJ517_ Net-_U6-PadJ518_ Net-_U6-PadJ519_ NC_19 MSP-EXP430F5529LP
U3 +3V3 Net-_U3-Pad2_ Net-_U3-Pad3_ NC_20 NC_21 NC_22 NC_23 NC_24 Net-_U3-Pad9_ GND NC_25 Net-_U3-Pad12_ Net-_U3-Pad13_ NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 XBee
U8 NC_33 Net-_U6-PadJ516_ Net-_U6-PadJ517_ Net-_U6-PadJ513_ Net-_U6-PadJ5.2_ Net-_U6-PadJ113_ NC_34 NC_35 Net-_U6-PadJ512_ Net-_U6-PadJ519_ NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 Net-_U6-PadJ5.4_ Net-_U6-PadJ518_ NC_43 NC_44 NC_45 Net-_U6-PadJ5.3_ Net-_U6-PadJ5.1_ OV7670
U7 NC_46 NC_47 NC_48 Net-_U6-PadJ517_ NC_49 Net-_U6-PadJ516_ NC_50 NC_51 NC_52 NC_53 Net-_U6-PadJ1.8_ NC_54 NC_55 NC_56 NC_57 NC_58 LPS331AP
U4 NC_59 GP-20U7
BT2 ~ GND Battery
BT1 NC_60 GND Battery
U2 ~ 3.6V
U1 ~ 3.6V
Q1 NC_61 Net-_Q1-Pad2_ NC_62 BUZ11
U5 ~ 3.6V
R1 ~ +3V3 R
R2 +3V3 GND R
Q2 Net-_Q2-Pad1_ Net-_Q2-Pad2_ +3V3 MMBT3904
Q3 Net-_Q3-Pad1_ Net-_Q3-Pad2_ +3V3 MMBT3904
R5 Net-_R5-Pad1_ GND R
TH1 Net-_Q2-Pad2_ Net-_R5-Pad1_ THERMISTOR
R6 Net-_Q3-Pad2_ Net-_R5-Pad1_ Photores
R3 NC_63 NC_64 R
R4 NC_65 NC_66 R
.end
