.title KiCad schematic
K_7 col0 NC_01 KEYSW
K_8 col1 NC_02 KEYSW
K_9 col2 NC_03 KEYSW
K_0 col3 NC_04 KEYSW
K_MINUS1 col4 NC_05 KEYSW
K_EQUAL1 col5 NC_06 KEYSW
K_BACKSPACE1 col6 NC_07 KEYSW
K_DEL1 col7 NC_08 KEYSW
K_Y1 col0 NC_09 KEYSW
K_U1 col1 NC_10 KEYSW
K_I1 col2 NC_11 KEYSW
K_O1 col3 NC_12 KEYSW
K_P1 col4 NC_13 KEYSW
K_[1 col5 NC_14 KEYSW
K_]1 col6 NC_15 KEYSW
K_BSLSH1 col7 NC_16 KEYSW
K_HOME1 NC_17 NC_18 KEYSW
K_H1 col0 NC_19 KEYSW
K_J1 col1 NC_20 KEYSW
K_K1 col2 NC_21 KEYSW
K_L1 col3 NC_22 KEYSW
K_SEMIC1 col4 NC_23 KEYSW
K_QUOTE1 col5 NC_24 KEYSW
K_ENTER1 col6 NC_25 KEYSW
K_END1 col7 NC_26 KEYSW
K_B1 col0 NC_27 KEYSW
K_N1 col1 NC_28 KEYSW
K_M1 col2 NC_29 KEYSW
K_COMMA1 col3 NC_30 KEYSW
K_DOT1 col4 NC_31 KEYSW
K_SLASH1 col5 NC_32 KEYSW
K_SHIFT1 col6 NC_33 KEYSW
K_5 col7 NC_34 KEYSW
K_`1 NC_35 NC_36 KEYSW
K_FN1 col0 NC_37 KEYSW
K_1 col1 NC_38 KEYSW
K_ALT1 col2 NC_39 KEYSW
K_CTRL1 col3 NC_40 KEYSW
K_2 col4 NC_41 KEYSW
K_3 col5 NC_42 KEYSW
K_4 col6 NC_43 KEYSW
.end
