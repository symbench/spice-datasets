.title KiCad schematic
R1 Net-_D1-Pad1_ Net-_C1-Pad1_ 470R
R2 Net-_BT1-Pad1_ Net-_C1-Pad2_ 47K
R4 Net-_D2-Pad1_ Net-_C2-Pad1_ 470R
R3 Net-_BT1-Pad1_ Net-_C2-Pad1_ 47K
D1 Net-_D1-Pad1_ Net-_BT1-Pad1_ LED
D2 Net-_D2-Pad1_ Net-_BT1-Pad1_ LED
BT1 Net-_BT1-Pad1_ Net-_BT1-Pad2_ 9V
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 47uF
C2 Net-_C2-Pad1_ Net-_C2-Pad1_ 47uF
U1 Net-_BT1-Pad2_ Net-_C2-Pad1_ Net-_C2-Pad1_ Net-_BT1-Pad2_ Net-_C1-Pad2_ Net-_C1-Pad1_ BC847RM
.end
