.title KiCad schematic
IC4 3.3VMCU NC_01 3.3VMCU 3.3VMCU NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 3.3VMCU NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 3.3VMCU NC_33 SCL NC_34 NC_35 SDA 3.3VMCU NC_36 NC_37 3.3VMCU NC_38 NC_39 NC_40 ESP32-PICO-D4
ANT1 NC_41 NC_42 NC_43 NC_44 ANT016008LCS2442MA1
AC1 NC_45 SDA NC_46 NC_47 NC_48 3.3VMCU 3.3VMCU NC_49 3.3VMCU SCL MC3635
.end
