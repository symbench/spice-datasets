.title KiCad schematic
SW1 Net-_D1-Pad1_ Net-_D2-Pad1_ Net-_D3-Pad1_ Earth Earth Earth SW_DIP_x03
D1 Net-_D1-Pad1_ Net-_D1-Pad2_ D
D2 Net-_D2-Pad1_ Net-_D2-Pad2_ D
D3 Net-_D3-Pad1_ Net-_D3-Pad2_ D
J1 Net-_D3-Pad2_ Net-_D2-Pad2_ Net-_D1-Pad2_ Conn_01x03
SW2 Net-_D4-Pad1_ Net-_D5-Pad1_ Net-_D6-Pad1_ Earth Earth Earth SW_DIP_x03
D4 Net-_D4-Pad1_ Net-_D4-Pad2_ D
D5 Net-_D5-Pad1_ Net-_D5-Pad2_ D
D6 Net-_D6-Pad1_ Net-_D6-Pad2_ D
J2 Net-_D6-Pad2_ Net-_D5-Pad2_ Net-_D4-Pad2_ Conn_01x03
SW3 Net-_D7-Pad1_ Net-_D8-Pad1_ Net-_D9-Pad1_ Earth Earth Earth SW_DIP_x03
D7 Net-_D7-Pad1_ Net-_D7-Pad2_ D
D8 Net-_D8-Pad1_ Net-_D8-Pad2_ D
D9 Net-_D9-Pad1_ Net-_D9-Pad2_ D
J3 Net-_D9-Pad2_ Net-_D8-Pad2_ Net-_D7-Pad2_ Conn_01x03
.end
