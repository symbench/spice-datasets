.title KiCad schematic
.include "/home/akshay/kicad-source-mirror-master/demos/simulation/sallen_key/ad8051.lib"
R3 Net-_C2-Pad1_ Net-_C1-Pad1_ 1k
R1 Net-_C1-Pad1_ ip 1k
R2 Net-_R2-Pad1_ GND 1k
R4 Net-_C1-Pad2_ Net-_R2-Pad1_ 1k
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 0.1u
C2 Net-_C2-Pad1_ GND 0.1u
V1 ip GND ac 1 0
R6 Net-_C3-Pad1_ Net-_C1-Pad2_ 1k
R7 Net-_C4-Pad1_ Net-_C3-Pad1_ 1k
C3 Net-_C3-Pad1_ out 0.1u
C4 Net-_C4-Pad1_ GND 0.1u
R5 Net-_R5-Pad1_ GND 1k
R8 out Net-_R5-Pad1_ 1k
V2 VDD GND dc 15
V3 GND VSS dc 15
XU1 Net-_R2-Pad1_ Net-_C2-Pad1_ VDD VSS Net-_C1-Pad2_ AD8051
XU2 Net-_R5-Pad1_ Net-_C4-Pad1_ VDD VSS out AD8051
.ac dec 10 1 1meg
.end
