.title KiCad schematic
R3 Net-_C3-Pad1_ /CANH0 60R
C3 Net-_C3-Pad1_ GND 47n
R1 Net-_C3-Pad1_ /CANL0 60R
C5 +3V3 GND 0.1u
C6 +3V3 GND 0.1u
C2 +3V3 GND 0.1u
C1 +3V3 GND 0.1u
IC1 +3V3 GND NC_01 NC_02 NC_03 NC_04 GND GND +3V3 GND NC_05 /CANH0 /CANL0 NC_06 GND GND ISO1050DW
IC2 +3V3 GND NC_07 NC_08 NC_09 NC_10 GND GND +3V3 GND NC_11 /CANH1 /CANL1 NC_12 GND GND ISO1050DW
R4 Net-_C4-Pad1_ /CANH1 60R
C4 Net-_C4-Pad1_ GND 47n
R2 Net-_C4-Pad1_ /CANL1 60R
.end
