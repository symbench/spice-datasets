.title KiCad schematic
D1 GND Net-_C1-Pad1_ Net-_C2-Pad2_ +3V3 PRTR5V0U2X
J1 NC_01 Net-_C1-Pad1_ Net-_C2-Pad2_ GND 5787834-1
R2 Net-_C2-Pad2_ NC_02 R
R1 Net-_C1-Pad1_ NC_03 R
C1 Net-_C1-Pad1_ GND C
C2 GND Net-_C2-Pad2_ C
J2 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 JD2-0001NL
IC1 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 NC_43 NC_44 NC_45 NC_46 NC_47 NC_48 NC_49 NC_50 NC_51 NC_52 NC_53 NC_54 NC_55 NC_56 NC_57 NC_58 NC_59 NC_60 NC_61 NC_62 NC_63 W5500
.end
