.title KiCad schematic
J1 /USB_1_SUPPLY Net-_J1-Pad2_ Net-_J1-Pad3_ GND GND USB_A
U2 Net-_J1-Pad3_ GND Net-_J2-Pad3_ Net-_J2-Pad2_ /5VIN Net-_J1-Pad2_ TPS2513A
U1 GND /5VIN /5VIN /~FAULT1 /~FAULT2 /~FAULT1 Net-_R3-Pad1_ /USB_2_SUPPLY /USB_1_SUPPLY /~FAULT2 GND TPS2561A
J2 /USB_2_SUPPLY Net-_J2-Pad2_ Net-_J2-Pad3_ GND GND USB_A
C5 /USB_1_SUPPLY GND CP1
C4 /USB_2_SUPPLY GND CP1
R3 Net-_R3-Pad1_ GND 25.5K
C1 /5VIN GND C
R1 /5VIN /~FAULT1 R
R2 /5VIN /~FAULT2 R
C2 /~FAULT1 GND 0.22uF
C3 /~FAULT2 GND 0.22uF
.end
