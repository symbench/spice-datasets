.title KiCad schematic
J1 /220_AC_Input/GND_in /220_AC_Input/220VAC 220VAC
J2 NC_01 /5V NC_02 /12V GNDREF Conn_01x05
T1 /220_AC_Input/220VAC /220_AC_Input/GND_in Net-_D1-Pad4_ Net-_D1-Pad3_ Transformer_1P_1S
D1 /12V/24V GNDREF Net-_D1-Pad3_ Net-_D1-Pad4_ D_Bridge_+-AA
C1 /12V/24V GNDREF 1500uF
U1 GNDREF /3.3V/3,3V /5V LM1117-3.3
C2 /5V GNDREF 10uF
C4 /3.3V/3,3V GNDREF 0,1uF
C3 /3.3V/3,3V GNDREF 22uF
U2 /12V /5V/GND /5V LM7805_TO220
C6 /5V /5V/GND C
C5 /12V /5V/GND C
U3 /12V GNDREF /9V/9V LM7809
C7 /12V GNDREF 0,1uF
C8 /9V/9V GNDREF 0,1uF
U4 /12V/24V GNDREF /12V LM7812
C9 /12V/24V GNDREF 0,1uF
C10 /12V GNDREF 0,1uF
.end
