.title KiCad schematic
U2 GND 32 33 25 26 27 DIO5 GND Net-_J7-Pad1_ GND DIO3 DIO4 +3V3 DIO0 DIO1 DIO2 RFM95HW
U1 GND +3V3 RESET NC_01 NC_02 34 35 32 33 25 26 27 14/SCL 12/SDA GND 13 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 15 2 0 4 16 17 5 18 19 NC_09 21 RX0 TX0 22 23/SAT_SLEEP GND GND ESP32-WROOM
J1 Net-_C1-Pad1_ GND +3V3 REG:3V3
C1 Net-_C1-Pad1_ GND 10 uF
C2 GND +3V3 22 uF
Q1 0 Net-_Q1-Pad2_ DTR Q_NPN_CBE
R2 Net-_Q1-Pad2_ RTS 10K
Q2 RESET Net-_Q2-Pad2_ RTS Q_NPN_CBE
R3 Net-_Q2-Pad2_ DTR 10K
J2 GND NC_10 VBUS RX0 TX0 RTS DTR prog
SW1 GND RESET SW_Push
R1 +3V3 RESET 10K
C3 RESET GND 1uF
SW2 GND 0 SW_Push
R4 +3V3 0 10K
C4 0 GND 1uF
J4 15 4 GND +3V3 16 GND 17 sdcard
J5 12/SDA 14/SCL GND +3V3 i2c-a
J7 Net-_J7-Pad1_ ANT
J8 +3V3 GND 12/SDA 14/SCL i2c-c
J9 GND 22 +3V3 1wire
J12 +3V3 18 NC_11 GND dht22
R7 +3V3 18 4.7K
J3 VIN GND VINS
R5 +3V3 12/SDA 4.7K
R6 +3V3 14/SCL 4.7K
J6 VIN GND +5V REG:5V
C5 VIN GND 10 uF
C6 GND +5V 22 uF
J14 SAT_RING_INDICATOR SAT_NETWORK_AVAIL 23/SAT_SLEEP SAT_LION satx
J15 +5V 35 21 19 5 2 0 VIN GND +3V3 14/SCL 12/SDA misc
J11 +3V3 VIN 21 19 GND uart
J19 GND +5V NC_12 SAT_RING_INDICATOR SAT_NETWORK_AVAIL 23/SAT_SLEEP SAT_LION GND 9602-b
J13 NC_13 34 13 +5V NC_14 GND 9602-a
R8 +3V3 22 R
J10 DIO2 DIO1 DIO0 +3V3 DIO4 DIO3 LBD
J16 33 32 26 25 DIO5 27 LBO
D1 Net-_C1-Pad1_ VBUS D
D2 Net-_C1-Pad1_ VIN D
.end
