.title KiCad schematic
J1 Net-_J1-Pad1_ GND Power conn
R2 Net-_R2-Pad1_ /in1 220
U2 Net-_R2-Pad1_ GNDD NC_01 GND Net-_R3-Pad1_ NC_02 4N35
R3 Net-_R3-Pad1_ VCC 10K
R4 Net-_R4-Pad1_ VCC 10K
R5 GND Net-_R4-Pad1_ 10K
Q1 VCC Net-_Q1-Pad2_ Net-_D2-Pad1_ BC547
Q2 GND Net-_Q1-Pad2_ Net-_D2-Pad1_ BC557
Q4 Net-_C6-Pad1_ Net-_J3-Pad2_ GND IRF3205
Q3 Net-_C6-Pad1_ Net-_J3-Pad2_ VCC IRF4905
R6 Net-_D2-Pad1_ Net-_C6-Pad1_ 10
D2 Net-_D2-Pad1_ Net-_C6-Pad1_ 1N4148
J3 Net-_J3-Pad1_ Net-_J3-Pad2_ MOTOR
J2 GNDD /in2 /in1 Input conn
R1 VCC Net-_D1-Pad2_ 5k
D1 GND Net-_D1-Pad2_ LED
U1 Net-_Q1-Pad2_ Net-_R3-Pad1_ Net-_R4-Pad1_ GND Net-_R8-Pad1_ Net-_R10-Pad1_ Net-_Q7-Pad2_ VCC LM358
R11 Net-_R11-Pad1_ /in2 220
U3 Net-_R11-Pad1_ GNDD NC_03 GND Net-_R10-Pad1_ NC_04 4N35
R10 Net-_R10-Pad1_ VCC 10k
R8 Net-_R8-Pad1_ VCC 10K
R9 GND Net-_R8-Pad1_ 10K
Q7 VCC Net-_Q7-Pad2_ Net-_D3-Pad1_ BC547
Q8 GND Net-_Q7-Pad2_ Net-_D3-Pad1_ BC557
Q6 Net-_C5-Pad1_ Net-_J3-Pad1_ GND IRF3205
Q5 Net-_C5-Pad1_ Net-_J3-Pad1_ VCC IRF4905
R7 Net-_D3-Pad1_ Net-_C5-Pad1_ 10
D3 Net-_D3-Pad1_ Net-_C5-Pad1_ 1N4148
C3 VCC GND C_Small
C4 VCC GND C_Small
C1 VCC GND CP
C2 VCC GND CP
J5 GNDD /in2 /in1 Input conn
J4 GNDD /in2 /in1 Input conn
C5 Net-_C5-Pad1_ VCC C_Small
C6 Net-_C6-Pad1_ VCC C_Small
SW1 Net-_J1-Pad1_ Net-_J1-Pad1_ VCC SW_SPDT
R12 Net-_D4-Pad2_ Net-_J1-Pad1_ 5k
D4 GND Net-_D4-Pad2_ LED
.end
