.title KiCad schematic
U3 +5V GND /SCL /SDA NC_01 /Temp NC_02 NC_03 Net-_D1-Pad2_ Net-_R1-Pad1_ /RES /SCK /MISO /MOSI /NSS +3V3 WeMos_mini
U1 +5V GND /SCL /SDA NC_04 NC_05 NC_06 NC_07 GY-521
R2 +3V3 /Temp 4.7k
R1 Net-_R1-Pad1_ +5V 220K
U5 GND /Temp +5V DS18B20
U4 NC_08 GND Net-_SW1-Pad1_ NC_09 NC_10 NC_11 TP4056-shield-6PIN
D1 /RES Net-_D1-Pad2_ Schottky
U2 GND GND +3V3 /RES NC_12 NC_13 NC_14 NC_15 GND NC_16 NC_17 /SCK /MISO /MOSI /NSS GND LoRa_Ra-02
SW2 Net-_SW1-Pad1_ +5V NC_18 SW_SPDT
SW1 Net-_SW1-Pad1_ +5V NC_19 SW_SPDT
C1 +5V GND 100n
.end
