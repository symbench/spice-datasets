.title KiCad schematic
U1 A14 A12 A7 A6 A5 A4 A3 A2 A1 A0 D0 D1 D2 NC_01 D3 D4 D5 D6 D7 NC_02 A10 ~RD A11 A9 A8 A13 NC_03 NC_04 LY62256PL-55LLI
U2 A14 A12 A7 A6 A5 A4 A3 A2 A1 A0 D0 D1 D2 NC_05 D3 D4 D5 D6 D7 NC_06 A10 ~RD A11 A9 A8 A13 NC_07 NC_08 LY62256PL-55LLI
.end
