.title KiCad schematic
R4 Net-_C1-Pad1_ 0 R
R2 Net-_R1-Pad2_ 0 R
R5 Net-_C3-Pad1_ 0 R
R3 +VDC Net-_C2-Pad1_ R
R1 +VDC Net-_R1-Pad2_ R
C5 Net-_C5-Pad1_ Net-_C4-Pad1_ C
C3 Net-_C3-Pad1_ Net-_C2-Pad1_ C
C4 Net-_C4-Pad1_ Net-_C3-Pad1_ C
C2 Net-_C2-Pad1_ NC_01 C
C1 Net-_C1-Pad1_ 0 C
Q1 Net-_C2-Pad1_ Net-_Q1-Pad2_ Net-_C1-Pad1_ NC_02 QNPN
R6 Net-_C4-Pad1_ 0 R
R7 Net-_C5-Pad1_ Net-_Q1-Pad2_ R_Variable
.end
