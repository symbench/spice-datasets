.title KiCad schematic
U1 NC_01 NC_02 GND +5V GND +5V NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 GND NC_17 Net-_R1-Pad1_ NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 ATmega328-AU
R1 Net-_R1-Pad1_ Net-_D1-Pad2_ R
D1 GND Net-_D1-Pad2_ LED
J1 GND +5V Conn_01x02_Female
.end
