.title KiCad schematic
TP1 NC_01 FID1
TP2 NC_02 FID1
.end
