.title KiCad schematic
J2 Net-_J1-Pad24_ Net-_J1-Pad23_ Net-_J1-Pad22_ Net-_J1-Pad21_ Net-_J1-Pad20_ Net-_J1-Pad19_ Net-_J1-Pad18_ Net-_J1-Pad17_ Net-_J1-Pad16_ Net-_J1-Pad15_ Net-_J1-Pad14_ Net-_J1-Pad13_ Net-_J1-Pad12_ Net-_J1-Pad11_ Net-_J1-Pad10_ Net-_J1-Pad9_ Net-_J1-Pad8_ Net-_J1-Pad7_ Net-_J1-Pad6_ Net-_J1-Pad5_ Net-_J1-Pad4_ Net-_J1-Pad3_ Net-_J1-Pad2_ Net-_J1-Pad1_ otp_FPC24
J1 Net-_J1-Pad1_ Net-_J1-Pad2_ Net-_J1-Pad3_ Net-_J1-Pad4_ Net-_J1-Pad5_ Net-_J1-Pad6_ Net-_J1-Pad7_ Net-_J1-Pad8_ Net-_J1-Pad9_ Net-_J1-Pad10_ Net-_J1-Pad11_ Net-_J1-Pad12_ Net-_J1-Pad13_ Net-_J1-Pad14_ Net-_J1-Pad15_ Net-_J1-Pad16_ Net-_J1-Pad17_ Net-_J1-Pad18_ Net-_J1-Pad19_ Net-_J1-Pad20_ Net-_J1-Pad21_ Net-_J1-Pad22_ Net-_J1-Pad23_ Net-_J1-Pad24_ Conn_01x24_Female
.end
