.title KiCad schematic
U1 Net-_J1-Pad6_ NC_01 NC_02 NC_03 NC_04 NC_05 +5V GNDPWR NC_06 NC_07 NC_08 NC_09 NC_10 Net-_R1-Pad1_ NC_11 NC_12 Net-_J1-Pad2_ Net-_J1-Pad10_ Net-_J1-Pad8_ +5V NC_13 GNDPWR NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 ATmega328-PU
J1 +5V Net-_J1-Pad2_ NC_20 NC_21 NC_22 Net-_J1-Pad6_ GNDPWR Net-_J1-Pad8_ NC_23 Net-_J1-Pad10_ SPI Connector
J2 +5V NC_24 GNDPWR NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 NC_43 GNDPWR Net-_J1-Pad8_ NC_44 Rainbow Bus
C1 +5V GNDPWR 100n
SW1 Net-_R1-Pad1_ +5V SW
R1 Net-_R1-Pad1_ GNDPWR 10k
D1 GNDPWR Net-_D1-Pad2_ LED_ALT
R2 Net-_D1-Pad2_ +5V 1k
C2 +5V GNDPWR 100u
.end
