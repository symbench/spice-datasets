.title KiCad schematic
R11 Net-_D7-Pad1_ Net-_P2-Pad6_ 1k
D7 Net-_D7-Pad1_ GND LED
D6 Net-_D6-Pad1_ GND LED
R10 Net-_D6-Pad1_ Net-_P2-Pad5_ 1k
R8 Net-_D4-Pad1_ Net-_P2-Pad3_ 1k
D4 Net-_D4-Pad1_ GND LED
D5 Net-_D5-Pad1_ GND LED
R9 Net-_D5-Pad1_ Net-_P2-Pad4_ 1k
R7 Net-_D3-Pad1_ Net-_P2-Pad2_ 1k
D3 Net-_D3-Pad1_ GND LED
D2 Net-_D2-Pad1_ GND LED
R6 Net-_D2-Pad1_ Net-_P2-Pad1_ 1k
K4 NC_01 COLONETTE
K2 NC_02 COLONETTE
K3 NC_03 COLONETTE
K1 NC_04 COLONETTE
C7 +5VD GND 47U
P3 GND Net-_P3-Pad2_ CONN_2
P8 Net-_P8-Pad1_ /SCL CAVALIER
P7 Net-_P7-Pad1_ /SDA CAVALIER
R5 Net-_P8-Pad1_ +5VD 2.1k
R4 Net-_P7-Pad1_ +5VD 2.1k
R3 /RST Net-_P3-Pad2_ 15
P6 GND /U2TX +5VD /U2RX CONN_4
D1 +5VD Net-_D1-Pad2_ LED
R2 Net-_D1-Pad2_ GND 1.5k
P2 Net-_P2-Pad1_ Net-_P2-Pad2_ Net-_P2-Pad3_ Net-_P2-Pad4_ Net-_P2-Pad5_ Net-_P2-Pad6_ CONN_6
C4 +5VD GND 6n8
C3 +5VD GND 6n8
C2 +5VD GND 6n8
C1 +5VD GND 6n8
SW1 GND Net-_P3-Pad2_ SW_PUSH_SMALL
C6 Net-_C6-Pad1_ GND 22p
C5 Net-_C5-Pad1_ GND 22p
X1 Net-_C5-Pad1_ Net-_C6-Pad1_ 7.3728Mhz
J1 /RST +5VD GND /PGD /PGC NC_05 NC_06 NC_07 RJ12
R1 +5VD Net-_P3-Pad2_ 10k
P4 GND +5VD /SCL /SDA CONN_4
P5 GND /U1ATX +5VD /U1ARX CONN_4
U1 Net-_P3-Pad2_ Net-_P2-Pad1_ Net-_P2-Pad2_ Net-_P2-Pad3_ Net-_P2-Pad4_ Net-_P2-Pad5_ Net-_P2-Pad6_ /PGC /PGD NC_08 +5VD GND Net-_C6-Pad1_ Net-_C5-Pad1_ /U1ATX /U1ARX NC_09 NC_10 NC_11 GND +5VD NC_12 NC_13 NC_14 /SCL /SDA /U2TX /U2RX NC_15 NC_16 GND +5VD NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 GND +5VD DSPIC30F4013
.end
