.title KiCad schematic
J1 BUS1 NC_01 BUS2 BUS20 BUS3 BUS21 BUS4 BUS22 BUS5 BUS23 BUS6 BUS24 BUS7 BUS25 BUS8 BUS26 BUS9 BUS27 BUS10 BUS28 BUS11 BUS29 BUS12 BUS30 BUS13 BUS31 BUS14 BUS32 BUS15 BUS33 BUS16 BUS34 BUS17 BUS35 BUS18 BUS36 BUS19 BUS37 NC_02 NC_03 PINS_2X20
U1 BUS1 BUS2 BUS3 BUS4 BUS5 BUS6 BUS7 BUS8 BUS9 BUS10 BUS11 BUS12 BUS13 BUS14 BUS15 BUS16 BUS17 BUS18 BUS19 BUS20 BUS21 BUS22 BUS23 BUS24 BUS25 BUS26 BUS27 BUS28 BUS29 BUS30 BUS31 BUS32 BUS33 BUS34 BUS35 BUS36 BUS37 BUS8 SUBD_2ROW_37PIN
U2 IFACE1 IFACE2 IFACE3 IFACE4 IFACE5 IFACE6 IFACE7 IFACE8 IFACE9 IFACE10 IFACE11 IFACE12 IFACE13 IFACE14 IFACE15 SUBD_2ROW_15PIN
J2 IFACE1 IFACE9 IFACE2 IFACE10 IFACE3 IFACE11 IFACE4 IFACE12 IFACE5 IFACE13 IFACE6 IFACE14 IFACE7 IFACE15 IFACE8 NC_04 PINS_2X08
.end
