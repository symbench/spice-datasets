.title KiCad schematic
SW2 GND NRST Reset
C4 +3V3 GND 4.7uF
C5 +3V3 GND 0.1uF
C6 +3V3 GND 0.1uF
C7 +3V3 GND 0.1uF
C8 +3V3 GND 0.1uF
C3 Net-_C3-Pad1_ GND 12pF
R4 Net-_C3-Pad1_ HSE_OUT 47
MH1 GND MountingHole_Pad
MH2 GND MountingHole_Pad
MH3 GND MountingHole_Pad
MH4 GND MountingHole_Pad
Y1 HSE_IN GND Net-_C3-Pad1_ GND Crystal_GND24
C1 HSE_IN GND 12pF
C2 NRST GND 0.1uF
J25 +3V3 SWDIO GND SWCLK GND SWO NC_01 NC_02 GND NRST SWD
C9 +3V3 GND 0.1uF
U1 +3V3 NC_03 NC_04 NC_05 HSE_IN HSE_OUT NRST NC_06 NC_07 NC_08 NC_09 GND +3V3 NC_10 NC_11 USART2_TX USART2_RX GND +3V3 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 USART3_TX USART3_RX GND +3V3 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 SWDIO GND +3V3 SWCLK NC_34 NC_35 NC_36 LCD_EN LCD_RS SWO LCD_D4 LCD_D5 I2C1_SCL I2C1_SDA GND LCD_D6 LCD_D7 GND +3V3 STM32F103RBT6
C11 GND +3V3 1uF
J27 +5V LCD_EN LCD_RS LCD_D4 LCD_D5 LCD_D6 LCD_D7 GND LCD
R2 +3V3 I2C1_SCL 4k7
R1 +3V3 I2C1_SDA 4k7
J29 +3V3 +3V3 +3V3 USART3_RX USART3_TX GND GND GND USART3
J28 +3V3 +3V3 +3V3 USART2_RX USART2_TX GND GND GND USART2
U3 GND +3V3 +5V AZ1117-3.3
C12 +5V GND 0.1uF
C13 +3V3 GND 0.1uF
J26 +5VP GND 5v In
D9 Net-_D9-Pad1_ +3V3 Power (Red)
R3 Net-_D9-Pad1_ GND 2k2
J30 +5VP +5VP +5V +5V 3557-2
.end
