.title KiCad schematic
U1 NC_01 GND NC_02 NC_03 GND NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 GND NC_12 NC_13 NC_14 Max4940
.end
