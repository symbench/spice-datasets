.title KiCad schematic
U1 NC_01 NC_02 Net-_U1-Pad14_ NC_03 NC_04 Net-_SW1-Pad1_ Net-_SW10-Pad1_ Net-_SW11-Pad1_ Net-_SW12-Pad1_ Net-_SW1-Pad2_ Net-_SW5-Pad2_ Net-_SW10-Pad2_ NC_05 Net-_U1-Pad14_ NC_06 NC_07 NC_08 NC_09 PIC_UNK
SW1 Net-_SW1-Pad1_ Net-_SW1-Pad2_ SWITCH_MOMENTARY
SW5 Net-_SW1-Pad1_ Net-_SW5-Pad2_ SWITCH_MOMENTARY
SW9 Net-_SW1-Pad1_ Net-_SW10-Pad2_ SWITCH_MOMENTARY
SW2 Net-_SW10-Pad1_ Net-_SW1-Pad2_ SWITCH_MOMENTARY
SW6 Net-_SW10-Pad1_ Net-_SW5-Pad2_ SWITCH_MOMENTARY
SW10 Net-_SW10-Pad1_ Net-_SW10-Pad2_ SWITCH_MOMENTARY
SW3 Net-_SW11-Pad1_ Net-_SW1-Pad2_ SWITCH_MOMENTARY
SW7 Net-_SW11-Pad1_ Net-_SW5-Pad2_ SWITCH_MOMENTARY
SW11 Net-_SW11-Pad1_ Net-_SW10-Pad2_ SWITCH_MOMENTARY
SW4 Net-_SW12-Pad1_ Net-_SW1-Pad2_ SWITCH_MOMENTARY
SW8 Net-_SW12-Pad1_ Net-_SW5-Pad2_ SWITCH_MOMENTARY
SW12 Net-_SW12-Pad1_ Net-_SW10-Pad2_ SWITCH_MOMENTARY
D4 NC_10 NC_11 LED_1206
D1 NC_12 Net-_D1-PadC_ LED_1206
D2 Net-_D1-PadC_ Net-_D2-PadC_ LED_1206
D3 Net-_D2-PadC_ NC_13 LED_1206
.end
