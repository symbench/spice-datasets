.title KiCad schematic
K1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 GND NC_07 FINDER-30.22
K2 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 GND NC_14 FINDER-30.22
K3 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 GND NC_21 FINDER-30.22
K4 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 GND NC_28 FINDER-30.22
.end
