.title KiCad schematic
V1 ip GND ac 5 0
R1 ip Net-_L1-Pad1_ 1k
L1 Net-_L1-Pad1_ GND 100m
C1 ip GND 0.1u
.ac dec 10 1 1meg
.end
