.title KiCad schematic
SD1 NC_01 SD_~CS SD_MOSI 3V3_PWR6 NC_02 GND SD_MISO NC_03 NC_04 NC_05 GND GND MICROSD
R23 SD_MISO 3V3_PWR6 47K
R24 SD_MOSI 3V3_PWR6 47K
R25 SD_~CS 3V3_PWR6 47K
.end
