.title KiCad schematic
J1 Net-_C1-Pad1_ Net-_J1-Pad2_ Net-_J1-Pad3_ Net-_J1-Pad4_ Net-_C1-Pad2_ Net-_C1-Pad2_ USB_B_Micro
J2 Net-_C1-Pad1_ Net-_J1-Pad2_ Net-_J1-Pad3_ Net-_J1-Pad4_ Net-_C1-Pad2_ USB
U1 Net-_C1-Pad2_ Net-_C2-Pad1_ Net-_C1-Pad1_ AMS1117-3.3
C2 Net-_C2-Pad1_ Net-_C1-Pad2_ 100n
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 100n
.end
