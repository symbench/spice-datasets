.title KiCad schematic
R201 NC_01 NC_02 1k
R202 NC_03 NC_04 1k
R203 NC_05 NC_06 1k
R204 NC_07 NC_08 1k
R205 NC_09 NC_10 1k
R206 NC_11 NC_12 1k
R207 NC_13 NC_14 1k
R208 NC_15 NC_16 1k
R301 NC_17 NC_18 1k
R302 NC_19 NC_20 1k
R303 NC_21 NC_22 1k
R304 NC_23 NC_24 1k
R305 NC_25 NC_26 1k
R306 NC_27 NC_28 1k
R307 NC_29 NC_30 1k
R308 NC_31 NC_32 1k
R401 NC_33 NC_34 1k
R402 NC_35 NC_36 1k
R403 NC_37 NC_38 1k
R404 NC_39 NC_40 1k
R405 NC_41 NC_42 1k
R406 NC_43 NC_44 1k
R407 NC_45 NC_46 1k
R408 NC_47 NC_48 1k
R501 NC_49 NC_50 1k
R502 NC_51 NC_52 1k
R503 NC_53 NC_54 1k
R504 NC_55 NC_56 1k
R505 NC_57 NC_58 1k
R506 NC_59 NC_60 1k
R507 NC_61 NC_62 1k
R508 NC_63 NC_64 1k
R601 NC_65 NC_66 1k
R602 NC_67 NC_68 1k
R603 NC_69 NC_70 1k
R604 NC_71 NC_72 1k
R605 NC_73 NC_74 1k
R606 NC_75 NC_76 1k
R607 NC_77 NC_78 1k
R608 NC_79 NC_80 1k
R701 NC_81 NC_82 1k
R702 NC_83 NC_84 1k
R703 NC_85 NC_86 1k
R704 NC_87 NC_88 1k
R705 NC_89 NC_90 1k
R706 NC_91 NC_92 1k
R707 NC_93 NC_94 1k
R708 NC_95 NC_96 1k
R801 NC_97 NC_98 1k
R802 NC_99 NC_100 1k
R803 NC_101 NC_102 1k
R804 NC_103 NC_104 1k
R805 NC_105 NC_106 1k
R806 NC_107 NC_108 1k
R807 NC_109 NC_110 1k
R808 NC_111 NC_112 1k
R901 NC_113 NC_114 1k
R902 NC_115 NC_116 1k
R903 NC_117 NC_118 1k
R904 NC_119 NC_120 1k
R905 NC_121 NC_122 1k
R906 NC_123 NC_124 1k
R907 NC_125 NC_126 1k
R908 NC_127 NC_128 1k
.end
