.title KiCad schematic
U1 GNDD /SPI_A0 /SPI_A1 /SPI_A2 NC_01 NC_02 NC_03 NC_04 NC_05 Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ Net-_U1-Pad16_ Net-_U1-Pad17_ /VIA_CLK /SPI5_MOSI +5V Net-_D1-Pad1_ NC_06 NC_07 +5V NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 W65C22S_PDIP
U3 +5V /SPI5_MISO Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ GNDD /SPI5_SCLK +5V Net-_U1-Pad14_ Net-_U1-Pad15_ Net-_U1-Pad16_ Net-_U1-Pad17_ +5V 74HC164
U2 GNDD /VIA_CLK NC_24 +5V NC_25 /SPI5_SCLK 74AC74
U604 /SPI_A0 /SPI_A1 /SPI_A2 GNDD GNDD +5V Net-_U604-Pad7_ GNDD Net-_U604-Pad9_ Net-_U604-Pad10_ Net-_U604-Pad11_ NC_26 NC_27 NC_28 NC_29 +5V 74HC138
D1 Net-_D1-Pad1_ NC_30 D
U605 NC_31 +3V3 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 Net-_R1-Pad2_ GNDD /SPI5_MOSI /SPI5_SCLK /SPI5_MISO NC_39 Net-_U604-Pad7_ Net-_U604-Pad9_ Net-_U604-Pad10_ +5V Net-_U604-Pad11_ TXS0108EPW
C1 +5V GNDD 100n
C2 +3V3 GNDD 100n
R1 /SPI_A2 Net-_R1-Pad2_ 2k7
R2 GNDD Net-_R1-Pad2_ 4k7
.end
