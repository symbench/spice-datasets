.title KiCad schematic
IC1 Net-_IC1-Pad1_ NC_01 NC_02 NC_03 NC_04 NC_05 Net-_IC1-Pad1_ LDL212PUR
IC2 Net-_IC2-Pad1_ NC_06 NC_07 NC_08 NC_09 NC_10 Net-_IC2-Pad1_ LDL212PUR
IC3 Net-_IC3-Pad1_ NC_11 NC_12 NC_13 NC_14 NC_15 Net-_IC3-Pad1_ LDL212PUR
.end
