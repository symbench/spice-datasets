.title KiCad schematic
P2 NC_01 +3V3 NC_02 +3V3 +5V GND GND NC_03 Power
P5 NC_04 NC_05 NC_06 GND NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 PWM
P3 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 Analog
P6 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 PWM
P4 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 Analog
P7 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 NC_43 NC_44 Communication
P1 GND GND NC_45 NC_46 NC_47 NC_48 NC_49 NC_50 NC_51 NC_52 NC_53 NC_54 NC_55 NC_56 NC_57 NC_58 NC_59 NC_60 NC_61 NC_62 NC_63 NC_64 NC_65 NC_66 NC_67 NC_68 NC_69 NC_70 NC_71 NC_72 NC_73 NC_74 NC_75 NC_76 +5V +5V Digital
Q2 NC_77 Earth Net-_J2-Pad1_ 2N7000
Ustep1 Net-_R[5v]1-Pad1_ NC_78 NC_79 NC_80 NC_81 NC_82 _
R[5v]1 Net-_R[5v]1-Pad1_ NC_83 R
J2 Net-_J2-Pad1_ CONN_01X01
J1 +5V CONN_01X01
Q3 NC_84 Earth Net-_J4-Pad1_ 2N7000
Udir1 Net-_R[5v]2-Pad1_ NC_85 NC_86 NC_87 NC_88 NC_89 _
R[5v]2 Net-_R[5v]2-Pad1_ NC_90 R
J4 Net-_J4-Pad1_ CONN_01X01
J3 +5V CONN_01X01
Q5 Net-_10K1-Pad2_ Earth Net-_J8-Pad1_ 2N7000
Uenab1 Net-_R[5v]4-Pad1_ NC_91 NC_92 NC_93 NC_94 NC_95 _
R[5v]4 Net-_R[5v]4-Pad1_ NC_96 R
J8 Net-_J8-Pad1_ CONN_01X01
J7 +5V CONN_01X01
Q1 NC_97 Earth Net-_10K1-Pad2_ 2N7000
10K1 +5V Net-_10K1-Pad2_ R
Q4 NC_98 Earth Net-_J6-Pad1_ 2N7000
Ustep2 Net-_R[5v]3-Pad1_ NC_99 NC_100 NC_101 NC_102 NC_103 _
R[5v]3 Net-_R[5v]3-Pad1_ NC_104 R
J6 Net-_J6-Pad1_ CONN_01X01
J5 +5V CONN_01X01
..../platform/atmel_sam/board/due/gShield-pinout.h 
.end
