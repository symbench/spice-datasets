.title KiCad schematic
D1 Net-_D1-Pad1_ Net-_D1-Pad2_ 0
R1 Net-_D1-Pad1_ Net-_R1-Pad2_ 1K
TP1 Net-_R1-Pad2_ 0
D2 Net-_D2-Pad1_ Net-_D1-Pad2_ 1
R2 Net-_D2-Pad1_ Net-_R2-Pad2_ 1K
TP2 Net-_R2-Pad2_ 1
D3 Net-_D3-Pad1_ Net-_D1-Pad2_ 2
R3 Net-_D3-Pad1_ Net-_R3-Pad2_ 1K
TP3 Net-_R3-Pad2_ 2
D4 Net-_D4-Pad1_ Net-_D1-Pad2_ 3
R4 Net-_D4-Pad1_ Net-_R4-Pad2_ 1K
TP4 Net-_R4-Pad2_ 3
D5 Net-_D5-Pad1_ Net-_D1-Pad2_ 4
R5 Net-_D5-Pad1_ Net-_R5-Pad2_ 1K
TP6 Net-_R5-Pad2_ 4
D6 Net-_D6-Pad1_ Net-_D1-Pad2_ 5
R6 Net-_D6-Pad1_ Net-_R6-Pad2_ 1K
TP7 Net-_R6-Pad2_ 5
D7 Net-_D7-Pad1_ Net-_D1-Pad2_ 6
R7 Net-_D7-Pad1_ Net-_R7-Pad2_ 1K
TP8 Net-_R7-Pad2_ 6
D8 Net-_D8-Pad1_ Net-_D1-Pad2_ 7
R8 Net-_D8-Pad1_ Net-_R8-Pad2_ 1K
TP9 Net-_R8-Pad2_ 7
TP5 Net-_D1-Pad2_ TEST
.end
