.title KiCad schematic
J11 Net-_J10-Pad1_ /D4- /D4+ Net-_J10-Pad4_ Net-_J10-Pad1_ /D3- /D3+ Net-_J10-Pad4_ Net-_J10-Pad4_ 2Port_USB2_0
J12 Net-_J10-Pad1_ /D7- /D7+ Net-_J10-Pad4_ Net-_J10-Pad1_ /D6- /D6+ Net-_J10-Pad4_ Net-_J10-Pad4_ 2Port_USB2_0
U3 /D4- /D4+ /D3- /D3+ D2- D2+ D1- D1+ NC_01 NC_02 NC_03 NC_04 /D6- /D6+ /D7- /D7+ Terminus_Technology_FE2.1
J10 Net-_J10-Pad1_ D1- D1+ Net-_J10-Pad4_ Net-_J10-Pad1_ D2- D2+ Net-_J10-Pad4_ Net-_J10-Pad4_ 2Port_USB2_0
.end
