.title KiCad schematic
U2 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 /QDR_D8 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 /QDR_D7 NC_43 NC_44 NC_45 NC_46 NC_47 NC_48 NC_49 NC_50 NC_51 /QDR_D6 NC_52 NC_53 NC_54 NC_55 NC_56 NC_57 NC_58 NC_59 NC_60 NC_61 NC_62 NC_63 NC_64 NC_65 NC_66 NC_67 NC_68 NC_69 NC_70 NC_71 NC_72 NC_73 /QDR_D5 NC_74 NC_75 NC_76 NC_77 NC_78 NC_79 NC_80 NC_81 NC_82 NC_83 NC_84 NC_85 NC_86 NC_87 NC_88 NC_89 NC_90 NC_91 NC_92 NC_93 NC_94 /QDR_D4 NC_95 NC_96 NC_97 NC_98 NC_99 NC_100 NC_101 NC_102 NC_103 /QDR_D3 NC_104 NC_105 NC_106 NC_107 NC_108 NC_109 NC_110 NC_111 NC_112 NC_113 NC_114 NC_115 NC_116 NC_117 NC_118 NC_119 NC_120 NC_121 NC_122 NC_123 NC_124 NC_125 /QDR_D2 NC_126 NC_127 NC_128 NC_129 NC_130 NC_131 NC_132 NC_133 NC_134 NC_135 /QDR_D1 NC_136 NC_137 NC_138 NC_139 NC_140 NC_141 NC_142 NC_143 NC_144 /QDR_D0 NC_145 NC_146 NC_147 NC_148 NC_149 NC_150 NC_151 NC_152 NC_153 NC_154 NC_155 NC_156 CY7C2245KV18-450BZKI
U1 NC_157 NC_158 NC_159 NC_160 NC_161 NC_162 NC_163 NC_164 NC_165 NC_166 NC_167 NC_168 NC_169 NC_170 NC_171 NC_172 NC_173 NC_174 NC_175 /QDR_D8 /QDR_D0 NC_176 NC_177 /QDR_D6 NC_178 NC_179 /QDR_D1 /QDR_D2 NC_180 NC_181 NC_182 /QDR_D7 NC_183 NC_184 /QDR_D3 NC_185 NC_186 NC_187 NC_188 NC_189 NC_190 /QDR_D4 /QDR_D5 NC_191 NC_192 NC_193 NC_194 NC_195 NC_196 NC_197 XC7KxT-FBG484
.end
