.title KiCad schematic
L6 +5V Net-_L6-Pad2_ GND Net-_L5-Pad2_ WS2812B
L1 +5V Net-_L1-Pad2_ GND Net-_L1-Pad4_ WS2812B
L20 +5V OUT_20Pixel GND Net-_L19-Pad2_ WS2812B
C19 +5V GND 104
C5 +5V GND 104
R1 Net-_L1-Pad4_ IN_20Pixel 471
P1 IN_20Pixel CONN_01X01
P2 GND CONN_01X01
P4 OUT_20Pixel CONN_01X01
P6 +5V CONN_01X01
P5 GND CONN_01X01
P3 +5V CONN_01X01
L2 +5V Net-_L2-Pad2_ GND Net-_L1-Pad2_ WS2812B
C1 +5V GND 104
L7 +5V Net-_L7-Pad2_ GND Net-_L6-Pad2_ WS2812B
C6 +5V GND 104
L12 +5V Net-_L12-Pad2_ GND Net-_L11-Pad2_ WS2812B
C11 +5V GND 104
L13 +5V Net-_L13-Pad2_ GND Net-_L12-Pad2_ WS2812B
C12 +5V GND 104
L14 +5V Net-_L14-Pad2_ GND Net-_L13-Pad2_ WS2812B
C13 +5V GND 104
L15 +5V Net-_L15-Pad2_ GND Net-_L14-Pad2_ WS2812B
C14 +5V GND 104
L16 +5V Net-_L16-Pad2_ GND Net-_L15-Pad2_ WS2812B
C15 +5V GND 104
L17 +5V Net-_L17-Pad2_ GND Net-_L16-Pad2_ WS2812B
C16 +5V GND 104
L18 +5V Net-_L18-Pad2_ GND Net-_L17-Pad2_ WS2812B
C17 +5V GND 104
L19 +5V Net-_L19-Pad2_ GND Net-_L18-Pad2_ WS2812B
C18 +5V GND 104
L3 +5V Net-_L3-Pad2_ GND Net-_L2-Pad2_ WS2812B
C2 +5V GND 104
L4 +5V Net-_L4-Pad2_ GND Net-_L3-Pad2_ WS2812B
C3 +5V GND 104
L5 +5V Net-_L5-Pad2_ GND Net-_L4-Pad2_ WS2812B
C4 +5V GND 104
L8 +5V Net-_L8-Pad2_ GND Net-_L7-Pad2_ WS2812B
C7 +5V GND 104
L9 +5V Net-_L10-Pad4_ GND Net-_L8-Pad2_ WS2812B
C8 +5V GND 104
L10 +5V Net-_L10-Pad2_ GND Net-_L10-Pad4_ WS2812B
C9 +5V GND 104
L11 +5V Net-_L11-Pad2_ GND Net-_L10-Pad2_ WS2812B
C10 +5V GND 104
.end
