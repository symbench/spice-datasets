.title KiCad schematic
.include "/home/akshay/Desktop/digital ciruits/libs/spice_models.lib"
X1 a b out VDD XOR
V1 a GND dc 0 pulse(0 3.3 0 0 0 50m 100m)
V3 VDD GND dc 3.3
V2 b GND dc 0 pulse(0 3.3 100m 0 0 50m 100m)
R1 GND out 10meg
.tran .25m 30m
.end
