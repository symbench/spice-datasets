.title KiCad schematic
U1 NC_01 GND NC_02 NC_03 NC_04 GND PYB30
.end
