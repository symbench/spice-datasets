.title KiCad schematic
MK1 NC_01 Mounting_Hole_PAD
MK2 NC_02 Mounting_Hole_PAD
MK3 NC_03 Mounting_Hole_PAD
MK4 NC_04 Mounting_Hole_PAD
.end
