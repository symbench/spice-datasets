.title KiCad schematic
IC1 /MOSI/SDA /MISO /SCK NC_01 VCC GND NC_02 NC_03 NC_04 /RESET NC_05 /RIGHT /ENC_A_RAW /ENC_B_RAW VCC GND /DOWN /OK /UP /LEFT TINY26S
R1 /RESET VCC 10k
R2 /ENC_B_RAW /ENC_B 10K
R3 /ENC_A_RAW /ENC_A 10K
C1 GND VCC 100n
C2 /ENC_A GND 100n
C3 /ENC_B GND 100n
BUTTONS1 /ENC_A /ENC_B GND GND /OK /DOWN /RIGHT /UP /LEFT ENCODER_ARROWS
POWER1 VCC NC_06 PINHD-1X2
OLED1 Net-_J2-Pad2_ Net-_J1-Pad2_ /SCK /MOSI/SDA PINHD-1X4
PROG1 /MOSI/SDA /MISO /SCK /RESET VCC GND PINHD-1X6
J1 GND Net-_J1-Pad2_ VCC SJ2W
J2 GND Net-_J2-Pad2_ VCC SJ2W
T1 NC_07 GND NC_08 AP2306GN_MOSFETSOT23
.end
