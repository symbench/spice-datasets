.title KiCad schematic
U1 +3V3 /P2 /P3 /P4 /P5 /P6 /P7 /P8 /P9 /P10 /P11 /P12 /P13 /P14 /P15 /~RST /TEST /P18 /P19 GND MSP430G2533IPW20
R1 Net-_D1-Pad1_ /P2 R_US
R3 +3V3 /~RST 47k
C4 /~RST GND 10nF
J1 +3V3 /P2 /P3 /P4 /P5 /P6 /P7 /P8 /P9 /P10 Conn_01x10
J2 /P11 /P12 /P13 /P14 /P15 /~RST /TEST /P18 /P19 GND Conn_01x10
D1 Net-_D1-Pad1_ +3V3 LED
R2 Net-_D2-Pad1_ GND R_US
D2 Net-_D2-Pad1_ +3V3 LED
C1 +3V3 GND 1uF
C2 +5V GND 10uF
C3 +3V3 GND 10uF
U2 GND +3V3 +5V AMS1117-3.3
J3 +5V NC_01 NC_02 NC_03 GND GND USB_B_Mini
SW1 GND /~RST SW_Push
.end
