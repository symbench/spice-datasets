.title KiCad schematic
U1 VCC_5V GND_BAT Net-_R1-Pad1_ 12V_DC/AC 12V_BAT ACS758
C2 GND_BAT IAC_DC C
C1 VCC_5V GND_BAT 0,1 uF
R1 Net-_R1-Pad1_ IAC_DC R
U2 VCC_5V GND_BAT Net-_R2-Pad1_ 12V_BAT +12V ACS758
C4 GND_BAT IBAT C
C3 VCC_5V GND_BAT 0,1 uF
R2 Net-_R2-Pad1_ IBAT R
U3 VCC_5V GND_BAT Net-_R3-Pad1_ 12V_Solarregler 12V_BAT ACS758
C6 GND_BAT I_Solarregler C
C5 VCC_5V GND_BAT 0,1 uF
R3 Net-_R3-Pad1_ I_Solarregler R
P1 VCC_5V IAC_DC GND_BAT IBAT NC_01 I_Solarregler NC_02 NC_03 12V_DC/AC NC_04 CONN_5X2
P2 12V_DC/AC CONN_1
P4 12V_BAT CONN_1
P3 12V_Solarregler CONN_1
.end
