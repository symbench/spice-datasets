.title KiCad schematic
P1 NC_01 NC_02 NC_03 +3V3 +5V GND GND NC_04 Power
P2 /A0 NC_05 NC_06 NC_07 /A4_SDA_ /A5_SCL_ Analog
P5 NC_08 CONN_01X01
P6 NC_09 CONN_01X01
P7 NC_10 CONN_01X01
P8 NC_11 CONN_01X01
P4 NC_12 NC_13 NC_14 GND NC_15 NC_16 NC_17 NC_18 Digital
P3 /A5_SCL_ /A4_SDA_ NC_19 GND NC_20 NC_21 NC_22 NC_23 NC_24 /8 Digital
D1 Net-_D1-Pad1_ /8 LED
RV1 +5V /A0 GND R_POT
SW1 +5V Net-_R1-Pad2_ SW_Push
R1 GND Net-_R1-Pad2_ R
R2 Net-_D1-Pad1_ GND R
.end
