.title KiCad schematic
J1 NC_01 NC_02 Net-_J1-Pad3_ NC_03 Net-_J1-Pad3_ NC_04 NC_05 NC_06 Net-_J1-Pad3_ NC_07 Conn_ARM_JTAG_SWD_10
.end
