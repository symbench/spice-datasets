.title KiCad schematic
U1 RPI_SEL NC_01 Net-_R5-Pad2_ NC_02 Net-_R6-Pad2_ NC_03 Net-_R7-Pad2_ NC_04 Net-_R8-Pad2_ GND NC_05 Net-_R4-Pad2_ NC_06 Net-_R3-Pad2_ NC_07 Net-_R2-Pad2_ NC_08 Net-_R1-Pad2_ RPI_SEL Net-_C1-Pad1_ 74HC244
U2 RPI_SEL Net-_U2-Pad2_ Net-_U2-Pad2_ Net-_R17-Pad2_ GND Net-_C1-Pad1_ 74HC04
R1 RPI_19 Net-_R1-Pad2_ 39k
R2 RPI_18 Net-_R2-Pad2_ 39k
R3 RPI_17 Net-_R3-Pad2_ 39k
R4 RPI_16 Net-_R4-Pad2_ 39k
R5 RPI_15 Net-_R5-Pad2_ 39k
R6 RPI_14 Net-_R6-Pad2_ 39k
R7 RPI_13 Net-_R7-Pad2_ 39k
R8 RPI_12 Net-_R8-Pad2_ 39k
R9 GND RPI_12 56κ
R10 GND RPI_13 56κ
R11 GND RPI_14 56κ
R12 GND RPI_15 56κ
R13 GND RPI_16 56κ
R14 GND RPI_17 56κ
R15 GND RPI_18 56κ
R16 GND RPI_19 56κ
R17 RPI_10 Net-_R17-Pad2_ 39k
R18 RPI_10 GND 56κ
C2 Net-_C1-Pad1_ GND 100n
C1 Net-_C1-Pad1_ GND 100n
.end
