.title KiCad schematic
R4 /ALT50HZ 5V 10K
RV2 /50HZ Net-_R3-Pad2_ Net-_R3-Pad2_ 10K
RV1 Net-_C1-Pad1_ Net-_R1-Pad1_ Net-_R1-Pad1_ 250K
R1 Net-_R1-Pad1_ Net-_C1-Pad1_ R
C1 Net-_C1-Pad1_ GND 100n
U2 GND Net-_C4-Pad1_ /50HZ 5V Net-_C2-Pad1_ Net-_C4-Pad1_ /ALT50HZ 5V TLC555
U1 GND /50HZ NC_01 5V Net-_C3-Pad1_ Net-_C1-Pad1_ Net-_C1-Pad1_ 5V TLC555
C3 Net-_C3-Pad1_ GND 100n
BT1 VIN GND Battery
P1 GND VIN CONN_01X02
C5 VIN GND 1U
R6 GND Net-_R5-Pad1_ R
R5 Net-_R5-Pad1_ 5V R
L1 VIN 5V INDUCTOR
U3 5V GND Net-_R5-Pad1_ VIN VIN AP3012
C6 5V GND C
C4 Net-_C4-Pad1_ GND .27U
C2 Net-_C2-Pad1_ GND 100n
R3 Net-_C4-Pad1_ Net-_R3-Pad2_ 46.4K
R2 5V Net-_R1-Pad1_ R
P2 GND VIN CONN_01X02
.end
