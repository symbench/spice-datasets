.title KiCad schematic
U1 GND +3V3 +5V +3V3 LM1117-3.3
C1 +3V3 GND CP
C2 +3V3 GND C
CON1 +5V GND MISO MOSI RXD SCK SCL SDA SSEL TXD UEXT-5V
J1 +3V3 +5V GND TXD RXD SCL SDA MISO MOSI SCK SSEL CONN_01X11
C3 +5V GND CP
CON2 +5V GND Net-_CON2-PadMISO_ Net-_CON2-PadMOSI_ Net-_CON2-PadRXD_ Net-_CON2-PadSCK_ Net-_CON2-PadSCL_ Net-_CON2-PadSDA_ Net-_CON2-PadSSEL_ Net-_CON2-PadTXD_ UEXT-BREADBOARD
CON3 +5V GND Net-_CON2-PadMISO_ Net-_CON2-PadMOSI_ Net-_CON2-PadRXD_ Net-_CON2-PadSCK_ Net-_CON2-PadSCL_ Net-_CON2-PadSDA_ Net-_CON2-PadSSEL_ Net-_CON2-PadTXD_ UEXT-5V
.end
