.title KiCad schematic
U5 NC_01 Net-_U5-Pad12_ Net-_U5-Pad10_ NC_02 NC_03 Net-_U5-Pad18_ Net-_U5-Pad18_ NC_04 NC_05 Net-_U5-Pad10_ NC_06 Net-_U5-Pad12_ NC_07 NC_08 NC_09 NC_10 Net-_U5-Pad17_ Net-_U5-Pad18_ Net-_U5-Pad18_ Net-_U5-Pad17_ NC_11 NC_12 NC_13 NC_14 L6235D
Alim12 NC_15 NC_16 B_Plug_5mm
.end
