.title KiCad schematic
J1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 +3V3 +3V3 GND NC_25 GND GND NC_26 VBAT VIN TEENSY3.2-72MHz
.end
