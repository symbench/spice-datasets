.title KiCad schematic
U2 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 BME680
U3 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 AS3935
R1 NC_25 NC_26 ALS-PT19-315C_L177_TR8
.end
