.title KiCad schematic
SW1 GND Net-_R1-Pad2_ RESET
SW2 Net-_R2-Pad1_ VCC INPUT_5
R2 Net-_R2-Pad1_ GND 10K
R3 SPKR+ PIN_6 220
R1 VCC Net-_R1-Pad2_ 10K
U1 PIN_1 Net-_R1-Pad2_ Net-_R2-Pad1_ GND PIN_5 PIN_6 PIN_7 VCC ATTINY85-20SU
J1 PIN_1 PIN_7 PIN_5 PIN_6 SPKR+ GND VCC GND Conn_01x08_Female
.end
