.title KiCad schematic
R2 Net-_C1-Pad1_ Net-_C1-Pad2_ 22
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 100p
C5 Net-_C1-Pad2_ Net-_C5-Pad2_ 220p
D1 Net-_D1-Pad1_ Net-_C1-Pad1_ BAT48 0.6V
D3 Net-_D3-Pad1_ Net-_C5-Pad2_ D1N4148
R6 Net-_C5-Pad2_ Net-_D3-Pad1_ 100k
R1 Net-_D3-Pad1_ Net-_D1-Pad1_ 1k
Q1 Net-_P1-Pad1_ Net-_C1-Pad1_ Net-_D1-Pad1_ Q2N2222
Q2 Net-_D3-Pad1_ Net-_C5-Pad2_ Net-_D1-Pad1_ Q2N2907
Q4 Net-_Q3-Pad1_ Net-_D1-Pad1_ Net-_P1-Pad1_ Q2N2907
Q6 Net-_C2-Pad2_ Net-_Q3-Pad1_ Net-_P1-Pad1_ Q2N2907
Q3 Net-_Q3-Pad1_ Net-_D1-Pad1_ Net-_D3-Pad1_ Q2N2222
Q5 Net-_C2-Pad2_ Net-_Q3-Pad1_ Net-_D3-Pad1_ Q2N2222
C2 Net-_C2-Pad1_ Net-_C2-Pad2_ 100n
C4 Net-_C4-Pad1_ Net-_C2-Pad2_ 100n
D5 Net-_D5-Pad1_ Net-_C4-Pad1_ BZD23-18
D2 Net-_C2-Pad1_ OUTPUT BZD23-18
R5 Net-_D5-Pad1_ Net-_C4-Pad1_ 1M
R3 Net-_C2-Pad1_ OUTPUT 1M
Q7 Net-_C4-Pad1_ Net-_Q7-Pad2_ Net-_D5-Pad1_ IRF9610
Q8 Net-_C2-Pad1_ Net-_Q7-Pad2_ OUTPUT IRF610
P1 Net-_P1-Pad1_ NC_01 NC_02 NC_03 NC_04 Net-_D3-Pad1_ NC_05 NC_06 Net-_C1-Pad2_ NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 CONN_01X19
P3 Net-_D5-Pad1_ NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 CONN_01X19
U1 OUTPUT Net-_D5-Pad1_ SMA
P2 OUTPUT Net-_P1-Pad1_ CONN_01X02
.end
