.title KiCad schematic
U1002 NC_01 NC_02 NC_03 GNDD Net-_U1001-Pad20_ +5V NC_04 GNDD NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 +5V 74HC138
C1002 +5V GNDD 100n
C1001 +5V GNDD 100n
U1001 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 GNDD NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 Net-_U1001-Pad20_ NC_29 NC_30 NC_31 +5V BUSCON_PDIP
.end
