.title KiCad schematic
J1 /MCLR Net-_J1-Pad2_ GND /ICSPDAT /ICSPCLK NC_01 HEADER_1X6
R11 Net-_R11-Pad1_ /ICSPDAT RES_0603
R12 Net-_R12-Pad1_ /ICSPCLK RES_0603
R5 Net-_C2-Pad1_ +3V3 RES_0603
C1 GND +3V3 CAP_0603
C2 Net-_C2-Pad1_ GND CAP_0603
U3 +3V3 NC_02 NC_03 /MCLR NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 Net-_R12-Pad1_ Net-_R11-Pad1_ GND PIC16F1829_SOIC
D1 Net-_C2-Pad1_ /MCLR Schottky_SMA
R6 +3V3 Net-_J1-Pad2_ RES_0603
.end
