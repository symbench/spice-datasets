.title KiCad schematic
U1 GND TRIGGER OUT RESET Net-_C2-Pad1_ THRESHOLD DISCHARGE VCC LM555
J1 GND VCC PWR
J2 VCC OUT GND OUT
C3 VCC GND 100nF
C2 Net-_C2-Pad1_ GND 100nF
R3 RESET VCC 10K
C1 THRESHOLD GND C_Small
x1 THRESHOLD DISCHARGE R_Small
x2 THRESHOLD TRIGGER R_Small
x3 RESET GND R_Small
x4 DISCHARGE GND R_Small
x5 TRIGGER VCC R_Small
x6 DISCHARGE VCC R_Small
D1 Net-_D1-Pad1_ VCC LED
R1 OUT Net-_D1-Pad1_ R_Small
D2 GND Net-_D2-Pad2_ LED
R2 OUT Net-_D2-Pad2_ R_Small
.end
