.title KiCad schematic
U1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 +5V GND NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 SCK MOSI MISO NC_18 NC_19 NC_20 Net-_R1-Pad2_ NC_21 NC_22 NC_23 RESET +5V GND Net-_C2-Pad1_ Net-_C3-Pad1_ NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 NC_43 NC_44 NC_45 NC_46 NC_47 NC_48 NC_49 +5V GND NC_50 NC_51 NC_52 NC_53 NC_54 NC_55 NC_56 NC_57 NC_58 NC_59 NC_60 NC_61 NC_62 NC_63 NC_64 NC_65 NC_66 +5V GND NC_67 NC_68 NC_69 NC_70 NC_71 NC_72 NC_73 NC_74 NC_75 NC_76 +5V GND Net-_C9-Pad1_ NC_77 NC_78 NC_79 NC_80 NC_81 NC_82 ATMEGA2560-16AUR
Y1 Net-_C2-Pad1_ Net-_C3-Pad1_ Crystal
C2 Net-_C2-Pad1_ GND C
C3 Net-_C3-Pad1_ GND C
R1 Net-_D1-Pad2_ Net-_R1-Pad2_ R
D1 GND Net-_D1-Pad2_ LED
R2 +5V RESET R
C4 +5V GND C
C5 +5V GND C
C6 +5V GND C
C7 +5V GND C
C8 +5V GND C
C9 Net-_C9-Pad1_ GND C
C10 RESET GND C
D2 Net-_C9-Pad1_ GND LM4040DBZ-3
R3 +5V Net-_C9-Pad1_ R
J1 MISO +5V SCK MOSI RESET GND AVR-ISP-6
J2 DTR NC_83 NC_84 +5V GND GND FTDI_Header
C1 RESET DTR C
.end
