.title KiCad schematic
SW1 Net-_J1-Pad2_ Net-_J1-Pad1_ SW_Push
J1 Net-_J1-Pad1_ Net-_J1-Pad2_ Conn_01x02_Female
.end
