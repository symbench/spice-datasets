.title KiCad schematic
C5 NC_01 Net-_C5-Pad2_ C
C7 NC_02 Net-_C5-Pad2_ C
C6 Net-_C6-Pad1_ NC_03 C
C8 Net-_C6-Pad1_ NC_04 C
J4 Net-_C5-Pad2_ NC_05 Net-_J4-Pad3_ Net-_J4-Pad3_ NC_06 Net-_C6-Pad1_ InConnector
J5 NC_07 NC_08 Net-_J5-Pad3_ Net-_J5-Pad3_ NC_09 NC_10 OutConnector
U2 NC_11 Net-_R10-Pad1_ NC_12 NC_13 NC_14 Net-_J5-Pad3_ NC_15 NC_16 OPA333xxD
R10 Net-_R10-Pad1_ Net-_J5-Pad3_ R
R7 NC_17 Net-_R6-Pad2_ R
R8 Net-_R6-Pad2_ Net-_J5-Pad3_ R
R9 Net-_R6-Pad2_ Net-_R10-Pad1_ R
R6 Net-_J4-Pad3_ Net-_R6-Pad2_ R
C13 NC_18 Net-_C13-Pad2_ C
C15 NC_19 Net-_C13-Pad2_ C
C14 Net-_C14-Pad1_ NC_20 C
C16 Net-_C14-Pad1_ NC_21 C
J8 Net-_C13-Pad2_ NC_22 Net-_J8-Pad3_ Net-_J8-Pad3_ NC_23 Net-_C14-Pad1_ InConnector
J9 NC_24 NC_25 Net-_J9-Pad3_ Net-_J9-Pad3_ NC_26 NC_27 OutConnector
R15 Net-_R14-Pad2_ Net-_R13-Pad2_ R
R12 NC_28 Net-_R11-Pad2_ R
R13 Net-_R11-Pad2_ Net-_R13-Pad2_ R
R14 Net-_R11-Pad2_ Net-_R14-Pad2_ R
R11 Net-_J8-Pad3_ Net-_R11-Pad2_ R
U3 Net-_R13-Pad2_ Net-_R14-Pad2_ NC_29 NC_30 NC_31 Net-_R19-Pad2_ Net-_J9-Pad3_ NC_32 ADA4807-2ARM
R20 Net-_R19-Pad2_ Net-_J9-Pad3_ R
R17 NC_33 Net-_R16-Pad2_ R
R18 Net-_R16-Pad2_ Net-_J9-Pad3_ R
R19 Net-_R16-Pad2_ Net-_R19-Pad2_ R
R16 Net-_R13-Pad2_ Net-_R16-Pad2_ R
.end
