.title KiCad schematic
N2 V20171120
N1 OHWLOGO
J1 NC_01 GNDA NC_02 NC_03 GNDA NC_04 GNDA NC_05 GNDA NC_06 GNDA NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 GND PINS_3X32
.end
