.title KiCad schematic
U1 DRIVE BAT SENSE TIMER SHDN PAUSE PROG ARCT SEL2 SEL1 NTC CHEM ACP +5V CHRG GND GND LTC4060
P2 GND CHRG +5V ACP CHEM NTC SEL1 SEL2 CONN_01X08
P1 ARCT PROG PAUSE SHDN TIMER SENSE BAT DRIVE CONN_01X08
.end
