.title KiCad schematic
J1 /IO02 /NC2 /IO00 /TMS /IO04 /IO34 /TDI /IO33 /IO32 /IO35 /IO25 /SVN /IO27 /NC1 /TD0 /TCK /5V /3.3V /GND /IO05 /IO16 /IO23 /IO17 /IO19 /SDA /IO18 /SCL /IO26 /RXD /SVP /TXD /RST Conn_02x16_Odd_Even
J3 /5V NC_01 /GND NC_02 /3.3V /IO04 /IO19 /GND /RXD /IO00 /TXD /GND /IO25 /IO33 /IO32 /IO35 /IO34 /RST /SVN /SVP Conn_02x10_Odd_Even
J2 /IO02 /NC2 /IO00 /TMS /IO04 /IO34 /TDI /IO33 /IO32 /IO35 /IO25 /SVN /IO27 /NC1 /TD0 /TCK /5V /3.3V /GND /IO05 /IO16 /IO23 /IO17 /IO19 /SDA /IO18 /SCL /IO26 /RXD /SVP /TXD /RST Conn_02x16_Odd_Even
J4 /3.3V /SCL /SDA /5V /GND Conn_01x05
.end
