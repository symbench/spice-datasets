.title KiCad schematic
J1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 QGND NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 Net-_J1-Pad15_ Net-_J1-Pad15_ QGND NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 FPC24
.end
