.title KiCad schematic
U1 GND MENB SCL SDA NC_01 +3V3 GND VOUT C2 C1 VREF WE RE CE GND LMP91002
P2 CE RE WE VREF C1 C2 VOUT CONN_01X07
P1 GND +3V3 NC_02 SDA SCL MENB GND CONN_01X07
.end
