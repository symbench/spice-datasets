.title KiCad schematic
U1 +BATT GND STBY NC_01 VOUT BU33SD5WG-TR
P1 VOUT +BATT GND STBY CONN_01X04
.end
