.title KiCad schematic
U2 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 +5V GND NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 GND +5V NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 PIC18F452-IP
U3 NC_37 NC_38 NC_39 LM324
.end
