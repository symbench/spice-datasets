.title KiCad schematic
U1 /A23 /A22 /A15 /A14 /A13 /A12 /A11 /A10 /A9 /A8 /A19 /A20 /~WE /~RST /A21 /~WP /RY~BY /A18 /A17 /A7 /A6 /A5 /A4 /A3 /A2 /A1 NC_01 NC_02 VDD NC_03 /A0 /~CS GND /~OE /D0 /D8 /D1 /D9 /D2 /D10 /D3 /D11 VCC /D4 /D12 /D5 /D13 /D6 /D14 /D7 /D15 GND /~BYTE /A16 /A25 /A24 EN29GL256
J1 /A0 /A1 /A2 /A3 /A4 /A5 /A6 /A7 /A8 /A9 /A10 /A11 /A12 /A13 /A14 /A15 /A16 /A17 /A18 /A19 /A20 /A21 /A22 /A23 /A24 /A25 ADDR
J2 /D14 /D15 /D12 /D13 /D10 /D11 /D8 /D9 /D6 /D7 /D4 /D5 /D2 /D3 /D0 /D1 GND VCC VDD /~BYTE /~CS /~OE /~RST /~WE /RY~BY /~WP DAT
C1 VCC GND 100nF
C2 VDD GND 100nF
.end
