.title KiCad schematic
R2 Net-_R1-Pad1_ Net-_R2-Pad2_ 2k
R1 Net-_R1-Pad1_ GND 2k
R4 Net-_R3-Pad1_ Net-_R4-Pad2_ 2k
R6 Net-_R5-Pad1_ Net-_R6-Pad2_ 2k
R8 Net-_R10-Pad2_ Net-_R8-Pad2_ 2k
R9 Net-_R10-Pad2_ GND 2k
R3 Net-_R3-Pad1_ Net-_R1-Pad1_ 1k
R5 Net-_R5-Pad1_ Net-_R3-Pad1_ 1k
R7 Net-_R10-Pad2_ Net-_R5-Pad1_ 1k
V1 Net-_R2-Pad2_ GND dc 0
V2 Net-_R4-Pad2_ GND dc 0
V3 Net-_R6-Pad2_ GND dc 0
V4 Net-_R8-Pad2_ GND dc 5
U1 out Net-_R10-Pad2_ GND AD8620
V5 VDD GND dc 10
V6 GND VSS dc 10
R10 out Net-_R10-Pad2_ 2k
.tran .25m 30m
.end
