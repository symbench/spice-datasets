.title KiCad schematic
U23 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 Net-_U23-Pad14_ NC_11 NC_12 Net-_U23-Pad17_ Net-_U23-Pad14_ NC_13 NC_14 NC_15 Net-_U23-Pad17_ NC_16 NC_17 NC_18 NC_19 NC_20 Net-_U23-Pad29_ NC_21 NC_22 Net-_U23-Pad29_ Net-_U23-Pad14_ NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 Net-_U23-Pad14_ NC_39 NC_40 NC_41 NC_42 NC_43 NC_44 NC_45 NC_46 NC_47 NC_48 NC_49 NC_50 NC_51 NC_52 NC_53 Net-_U23-Pad17_ IDT7005J
.end
