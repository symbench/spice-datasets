.title KiCad schematic
U1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 74HC109
.end
