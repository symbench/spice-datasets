.title KiCad schematic
J2 Net-_J1-Pad16_ NC_01 GND NC_02 GND NC_03 GND NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 GND NC_11 GND GND GND NC_12 NC_13 NC_14 NC_15 GND ATX24
D1 NC_16 NC_17 LED
D2 NC_18 NC_19 LED
J1 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 Net-_J1-Pad16_ NC_35 NC_36 CONN_02X09
J3 Net-_J1-Pad16_ NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 NC_43 NC_44 NC_45 NC_46 NC_47 NC_48 NC_49 NC_50 NC_51 NC_52 NC_53 NC_54 NC_55 NC_56 NC_57 NC_58 NC_59 ATX_24PIN
.end
