.title KiCad schematic
N2 V20190807
N1 OHWLOGO
.end
