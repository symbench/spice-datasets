.title KiCad schematic
P3 NC_01 CONN_01X01
P4 NC_02 CONN_01X01
P5 NC_03 CONN_01X01
P6 NC_04 CONN_01X01
P1 NC_05 NC_06 /Reset GND NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 Digital
P2 NC_18 GND /Reset +5V NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 +3V3 NC_28 Analog
.end
