.title KiCad schematic
K1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 OMRON-G2R-24
.end
