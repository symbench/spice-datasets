.title KiCad schematic
U3 GND +3V3 /EN NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 GND NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 /IO2 /IO0 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 /RXD0 /TXD0 NC_28 NC_29 GND GND ESP32-WROOM-32
R3 +3V3 /EN 10kR
C1 /EN GND 0.1uF
C5 +3V3 GND 0.1uF
C4 +3V3 GND 22uF
C2 GND /IO0 0.1uF
SW2 GND /IO0 BOOT
C3 GND /EN 0.1uF
SW3 GND /EN RESET
J5 /RXD0 +3V3 /IO0 NC_30 /IO2 NC_31 GND /TXD0 Conn_02x04_Odd_Even
.end
