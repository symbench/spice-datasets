.title KiCad schematic
D1 Net-_C1-Pad1_ Net-_D1-Pad2_ 1N60
R1 NC_01 Net-_C1-Pad2_ 3.9k
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 10p
P1 Net-_C1-Pad2_ NC_02 NC_03 Net-_D1-Pad2_ NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 CONN_01X19
P2 NC_19 NC_20 NC_21 NC_22 Net-_C1-Pad1_ NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 CONN_01X19
.end
