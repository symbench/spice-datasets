.title KiCad schematic
R18 +3V3 SWCLK 1k
C29 RST GND 100nF
SW1 GND Net-_R17-Pad1_ RESET
R17 Net-_R17-Pad1_ RST 330
R15 +3V3 RST 10k
U5 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 GND +3V3 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 GND Net-_U5-Pad25_ FLASH_MOSI FLASH_SCK FLASH_CS FLASH_MISO Net-_U5-Pad25_ GND NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 GND +3V3 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 GND +3V3 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 NC_43 NC_44 NC_45 NC_46 GND +3V3 NC_47 NC_48 NC_49 NC_50 NC_51 NC_52 NC_53 NC_54 NC_55 NC_56 NC_57 NC_58 GND +3V3 NC_59 NC_60 NC_61 NC_62 NC_63 NC_64 NC_65 NC_66 NC_67 NC_68 RST VDDCORE GND VSW +3V3 SWCLK NC_69 NC_70 NC_71 NC_72 NC_73 NC_74 NC_75 SAMD51
R16 +3V3 FLASH_CS 10k
C21 +3V3 GND 10uF
C22 +3V3 GND 10uF
C23 +3V3 GND 10uF
C24 +3V3 GND 10uF
C25 +3V3 GND 10uF
C26 +3V3 GND 100nF
C27 VDDCORE GND 4.7uF
C28 VDDCORE GND 100nF
L2 VDDCORE VSW 10uH
U6 FLASH_CS FLASH_MISO FLASH_CS GND FLASH_MOSI FLASH_SCK FLASH_CS +3V3 AT25DF041B-SSHN-T
.end
