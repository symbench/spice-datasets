.title KiCad schematic
DS1 GND +5V Net-_DS1-Pad3_ Net-_DS1-Pad4_ GND Net-_DS1-Pad6_ NC_01 NC_02 NC_03 NC_04 Net-_DS1-Pad11_ Net-_DS1-Pad12_ Net-_DS1-Pad13_ Net-_DS1-Pad14_ Net-_DS1-Pad15_ GND WC1602A
U2 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 Net-_DS1-Pad14_ Net-_DS1-Pad13_ Net-_DS1-Pad12_ Net-_DS1-Pad11_ NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 Net-_DS1-Pad6_ Net-_DS1-Pad4_ NC_21 +3V3 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 Net-_U1-Pad2_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad3_ NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 STM32F103C8Tx
U1 GND Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ NC_42 GND +3V3 BME280
R220 +5V Net-_DS1-Pad15_ R
R_Poti1 GND Net-_DS1-Pad3_ +5V 10kOhm
.end
