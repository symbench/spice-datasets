.title KiCad schematic
U201 Net-_C504-Pad1_ PP_USB /USB2_DM /USB1_DM PP_USB /USB2_DP /USB1_DP NC_01 MCIMX6Y2DVM
C504 Net-_C504-Pad1_ COM 0.22u
C505 Net-_C504-Pad1_ COM 10u
C503 PP_USB COM 1u
C502 PP_USB COM 1u
J501 PP_USB_DEVICE /USB1_DM /USB1_DP NC_02 COM COM USB-MICROB
J502 /PP_USB_HOST /USB1_DP /USB1_DM COM COM USB-HEADER-5PIN
U501 PP_USB COM PP_USB /PP_USB_HOST /USB1_DM /USB1_DP TPD3S014
C507 /PP_USB_HOST COM 120u
C506 PP_USB COM 0.22u
R501 PP_USB /PP_USB_HOST 0
M501 PP_WLAN Net-_J503-Pad1_ COM /USB2_DM /USB2_DP RTL8188EUS
C508 PP_WLAN COM 22u
J503 Net-_J503-Pad1_ COM CONN-2
C501 PP_USB_DEVICE COM 10u
.end
