.title KiCad schematic
K1 Net-_J3-Pad2_ Net-_J3-Pad1_ Net-_J3-Pad3_ Net-_D1-Pad2_ Net-_D1-Pad1_ FINDER-40.31
J1 GND Net-_J1-Pad2_ VCC Conn_01x03
U1 Net-_R1-Pad1_ GND Net-_D1-Pad2_ Net-_R2-Pad2_ PC817
R1 Net-_R1-Pad1_ Net-_J1-Pad2_ 1k
JP2 GND Net-_D1-Pad2_ Jumper
JP1 VCC Net-_J4-Pad1_ Jumper
J3 Net-_J3-Pad1_ Net-_J3-Pad2_ Net-_J3-Pad3_ Conn_01x03
J4 Net-_J4-Pad1_ Conn_01x01
J2 Net-_D1-Pad2_ Conn_01x01
D1 Net-_D1-Pad1_ Net-_D1-Pad2_ D_Small
Q1 Net-_Q1-Pad1_ Net-_J4-Pad1_ Net-_D1-Pad1_ Q_PNP_BEC
R2 Net-_Q1-Pad1_ Net-_R2-Pad2_ 1k
R3 Net-_Q1-Pad1_ Net-_J4-Pad1_ 1k
.end
