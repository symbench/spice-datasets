.title KiCad schematic
K_ESC1 col0 NC_01 KEYSW
K_DEL1 col1 NC_02 KEYSW
K_1 col2 NC_03 KEYSW
K_2 col3 NC_04 KEYSW
K_3 col4 NC_05 KEYSW
K_4 col5 NC_06 KEYSW
K_5 col6 NC_07 KEYSW
K_6 NC_08 NC_09 KEYSW
K_END1 col0 NC_10 KEYSW
K_TAB1 col1 NC_11 KEYSW
K_Q1 col2 NC_12 KEYSW
K_W1 col3 NC_13 KEYSW
K_E1 col4 NC_14 KEYSW
K_R1 col5 NC_15 KEYSW
K_T1 col6 NC_16 KEYSW
K_HOME1 col0 NC_17 KEYSW
K_CAPS_LOCK1 col1 NC_18 KEYSW
K_A1 col2 NC_19 KEYSW
K_S1 col3 NC_20 KEYSW
K_D1 col4 NC_21 KEYSW
K_F1 col5 NC_22 KEYSW
K_G1 col6 NC_23 KEYSW
K_`1 col0 NC_24 KEYSW
K_SHIFT1 col1 NC_25 KEYSW
K_Z1 col2 NC_26 KEYSW
K_X1 col3 NC_27 KEYSW
K_C1 col4 NC_28 KEYSW
K_V1 col5 NC_29 KEYSW
K_FN1 col0 NC_30 KEYSW
K_CTRL1 col1 NC_31 KEYSW
K_ALT1 col2 NC_32 KEYSW
K_7 col3 NC_33 KEYSW
.end
