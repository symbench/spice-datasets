.title KiCad schematic
U2 Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U2-Pad7_ Net-_U2-Pad8_ Net-_U2-Pad9_ Net-_U2-Pad10_ Net-_U2-Pad11_ Net-_U2-Pad12_ Net-_U2-Pad13_ NC_01 Net-_U2-Pad15_ Net-_U2-Pad16_ Net-_U2-Pad17_ Net-_U2-Pad18_ Net-_U2-Pad19_ NC_02 Net-_U2-Pad21_ Net-_U2-Pad22_ Net-_U2-Pad23_ Net-_U2-Pad24_ Net-_U2-Pad25_ Net-_U2-Pad26_ NC_03 NC_04 LY62256PL-55LLI
U3 Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U2-Pad7_ Net-_U2-Pad8_ Net-_U2-Pad9_ Net-_U2-Pad10_ Net-_U2-Pad11_ Net-_U2-Pad12_ Net-_U2-Pad13_ NC_05 Net-_U2-Pad15_ Net-_U2-Pad16_ Net-_U2-Pad17_ Net-_U2-Pad18_ Net-_U2-Pad19_ NC_06 Net-_U2-Pad21_ Net-_U2-Pad22_ Net-_U2-Pad23_ Net-_U2-Pad24_ Net-_U2-Pad25_ Net-_U2-Pad26_ NC_07 NC_08 LY62256PL-55LLI
.end
