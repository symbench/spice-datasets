.title KiCad schematic
U1 VOUT_UC Net-_R2-Pad1_ Net-_R3-Pad2_ GND VCC LM358
R3 VCC Net-_R3-Pad2_ 10K
R4 Net-_R3-Pad2_ GND 10K
R5 VOUT_UC Net-_R2-Pad1_ 100K
R1 VCC MIC 10K
R2 Net-_R2-Pad1_ Net-_CP1-Pad2_ 1K
CP1 MIC Net-_CP1-Pad2_ 10uF
CP2 VOUT_UC VOUT 220uF
C1 VCC GND 100nF
P1 GND MIC CONN_01X02
P2 GND VOUT CONN_01X02
P3 GND VOUT_UC CONN_01X02
P4 GND VCC CONN_01X02
.end
