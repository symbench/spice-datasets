.title KiCad schematic
R1 +3V3 Temp_0 4K7
R2 +3V3 Temp_1 4k7
J2 +5V GND NC_01 Endstop_X
C2 Temp_1 GND 10uF
C1 Temp_0 GND 10uF
R5 GND Hotend 10k
R6 GND Heatbed 10k
J3 GND +5V Servo_0_Buff Servo_0
J1 +3V3 GND SDA SCL I2C
J7 +3V3 GND MISO_2 MOSI_2 SCK_2 SDCS SPI
J33 Temp_1 GND TEMP_1
J32 Temp_0 GND TEMP_0
J5 GND +5V Servo_1_Buff Servo_1
J4 +5V GND NC_02 Endstop_Y
J6 +5V GND NC_03 Endstop_Z
C3 +5V GND 100nF
J16 +3V3 +3V3 GND GND NC_04 NC_05 NC_06 NC_07 Serial_1_2
J27 +3V3 +3V3 GND GND NC_08 NC_09 PB12 PB13 Serial_3_4
D1 GND Net-_D1-Pad2_ LED_RED
R3 Net-_D1-Pad2_ PB12 150R
D2 GND Net-_D2-Pad2_ LED_RED
R4 Net-_D2-Pad2_ PB13 150R
J8 NC_10 Net-_J30-Pad5_ GND GPIO0_SEL
R26 +3V3 SCL 4k7
R27 +3V3 SDA 4k7
J29 NC_11 SDCS MOSI_2 +3V3 SCK_2 GND MISO_2 NC_12 NC_13 GND Micro_SD_Card_Det
U3 GND Heatbed NC_14 GND Hotend NC_15 GND Servo_1_Buff NC_16 GND Servo_0_Buff NC_17 GND +5V 74HCT125
J30 GND NC_18 NC_19 +3V3 Net-_J30-Pad5_ NC_20 NC_21 +3V3 ESP-01v090
.end
