.title KiCad schematic
C92 NC_01 Net-_C92-Pad2_ C
C94 NC_02 Net-_C92-Pad2_ C
C93 Net-_C93-Pad1_ NC_03 C
C95 Net-_C93-Pad1_ NC_04 C
J34 Net-_C92-Pad2_ NC_05 Net-_C96-Pad2_ Net-_C96-Pad2_ NC_06 Net-_C93-Pad1_ InConnector
J35 NC_07 NC_08 Net-_C97-Pad1_ Net-_C97-Pad1_ NC_09 NC_10 OutConnector
U20 NC_11 Net-_R240-Pad1_ Net-_C96-Pad1_ NC_12 NC_13 Net-_C97-Pad2_ NC_14 NC_15 OPA333xxD
R242 NC_16 Net-_C96-Pad1_ R
R241 Net-_C96-Pad2_ Net-_C97-Pad1_ R
R240 Net-_R240-Pad1_ Net-_C96-Pad2_ R
C97 Net-_C97-Pad1_ Net-_C97-Pad2_ C
C96 Net-_C96-Pad1_ Net-_C96-Pad2_ C
R243 Net-_R240-Pad1_ Net-_C97-Pad2_ R
.end
