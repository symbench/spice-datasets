.title KiCad schematic
J2 VBUS NC_01 NC_02 NC_03 GND GND USB_B_Micro
J1 NC_04 GND Jack-DC
U1 Net-_U1-Pad1_ NC_05 NC_06 Net-_U1-Pad4_ Net-_U1-Pad4_ NC_07 NC_08 Net-_U1-Pad1_ USB6B1
Y1 NC_09 NC_10 Crystal
U2 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 GND NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 GND NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 GND NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 GND NC_41 NC_42 NC_43 NC_44 NC_45 NC_46 NC_47 NC_48 NC_49 NC_50 GND NC_51 GND NC_52 FT2232D
.end
