.title KiCad schematic
U3 NC_01 /Diagnostic Net-_U3-Pad10_ NC_02 NC_03 Net-_U3-Pad18_ Net-_U3-Pad18_ NC_04 NC_05 Net-_U3-Pad10_ NC_06 /Diagnostic NC_07 NC_08 NC_09 NC_10 Net-_U3-Pad17_ Net-_U3-Pad18_ Net-_U3-Pad18_ Net-_U3-Pad17_ NC_11 NC_12 NC_13 NC_14 L6235PD
.end
