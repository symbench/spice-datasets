.title KiCad schematic
U8 /VIN_UNREG NC_01 NC_02 /VIN_UNREG NC_03 NC_04 TLV62568DDC
.end
