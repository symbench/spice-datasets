.title KiCad schematic
X1 Net-_C3-Pad1_ GND Net-_C4-Pad1_ GND 16MHz 18pF
C2 +12V GND 10uF 25V
C6 Net-_C6-Pad1_ GND 10uF 25V
C3 Net-_C3-Pad1_ GND 22pF
C4 Net-_C4-Pad1_ GND 22pF
D1 /VIN GND 14V
F1 +12V Net-_D2-Pad1_ 1.1A 25V
J1 /VIN GND INPUT
D2 Net-_D2-Pad1_ /VIN 20V 1A
C7 +5V GND 100nF
C8 +5V GND 100nF
C9 +5V GND 100nF
S1 GND /~RESET RESET
J3 /D11 +5V /D13 /D12 /~RESET GND ISP-2560
U1 GND Net-_C6-Pad1_ +12V NCP1117-5V
C1 /~RESET /FTDI_RESET 100nF
J2 /FTDI_RESET /D0 /D1 +5V NC_01 GND FTDI
D3 +5V Net-_C6-Pad1_ 20V 1A
LED1 GND NC_02 AMBER
C5 +5V GND 100nF
U2 /D3 /D4 GND +5V GND +5V Net-_C3-Pad1_ Net-_C4-Pad1_ /D5 /D6 /D7 /D8 /D9 /D10 /D12 /D11 /D13 +5V /A6_*_ +5V GND /A7_*_ /A0 /A1 /A2 /A3 /A4 /A5 /~RESET /D0 /D1 /D2 ATMEGA328
J4 /D2 /D3 /D4 /D5 /D6 /D7 /D8 /D9 /D10 /D11 DIGOUT1
J5 /D12 /D13 /A0 /A1 /A2 /A3 /A4 /A5 /A6_*_ /A7_*_ DIGOUT2
.end
