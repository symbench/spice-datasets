.title KiCad schematic
U9 3.3V 3.3V 3.3V GND NC_01 NC_02 GND 3.3V MB85RC256
.end
