.title KiCad schematic
J1 Net-_J1-Pad1_ Net-_J1-Pad2_ Net-_J1-Pad3_ NC_01 Net-_J1-Pad5_ Net-_J1-Pad5_ USB_B_Micro
J2 Net-_J1-Pad1_ Net-_J1-Pad2_ Net-_J1-Pad3_ NC_02 Net-_J1-Pad5_ Net-_J1-Pad5_ USB_B_Micro
.end
