.title KiCad schematic
U1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 +5V GND NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 GND +5V Net-_D1-Pad2_ Net-_D2-Pad2_ Net-_D3-Pad2_ Net-_D4-Pad2_ Net-_D5-Pad2_ Net-_D6-Pad2_ Net-_D7-Pad2_ Net-_D8-Pad2_ PIC18F4550-IP
D3 Net-_D3-Pad1_ Net-_D3-Pad2_ LED
D4 Net-_D4-Pad1_ Net-_D4-Pad2_ LED
D5 Net-_D5-Pad1_ Net-_D5-Pad2_ LED
D6 Net-_D6-Pad1_ Net-_D6-Pad2_ LED
D7 Net-_D7-Pad1_ Net-_D7-Pad2_ LED
D2 Net-_D2-Pad1_ Net-_D2-Pad2_ LED
D1 Net-_D1-Pad1_ Net-_D1-Pad2_ LED
D8 Net-_D8-Pad1_ Net-_D8-Pad2_ LED
R1 Net-_D1-Pad1_ GND R
R2 Net-_D2-Pad1_ GND R
R3 Net-_D3-Pad1_ GND R
R4 Net-_D4-Pad1_ GND R
R5 Net-_D5-Pad1_ GND R
R6 Net-_D6-Pad1_ GND R
R7 Net-_D7-Pad1_ GND R
R8 Net-_D8-Pad1_ GND R
.end
