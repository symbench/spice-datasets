.title KiCad schematic
U4 GND NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 VCC NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 GND GND NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 VCC NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 WD65C816S_PLCC44-65xx
C7 GND VCC 0.1uF
C6 VCC GND 0.1uF
U1 NC_40 NC_41 NC_42 NC_43 NC_44 NC_45 NC_46 NC_47 Net-_U1-Pad27_ Net-_U1-Pad10_ NC_48 NC_49 NC_50 NC_51 NC_52 NC_53 NC_54 NC_55 NC_56 NC_57 NC_58 NC_59 NC_60 NC_61 NC_62 NC_63 Net-_U1-Pad27_ Net-_U1-Pad10_ NC_64 NC_65 NC_66 NC_67 NC_68 NC_69 NC_70 NC_71 IS61C5128AL-10KLI
U2 NC_72 NC_73 NC_74 NC_75 NC_76 NC_77 NC_78 NC_79 Net-_U2-Pad27_ Net-_U2-Pad10_ NC_80 NC_81 NC_82 NC_83 NC_84 NC_85 NC_86 NC_87 NC_88 NC_89 NC_90 NC_91 NC_92 NC_93 NC_94 NC_95 Net-_U2-Pad27_ Net-_U2-Pad10_ NC_96 NC_97 NC_98 NC_99 NC_100 NC_101 NC_102 NC_103 IS61C5128AL-10KLI
U3 NC_104 NC_105 NC_106 NC_107 NC_108 NC_109 NC_110 NC_111 NC_112 NC_113 NC_114 NC_115 NC_116 NC_117 NC_118 NC_119 NC_120 NC_121 NC_122 NC_123 NC_124 NC_125 NC_126 NC_127 NC_128 NC_129 NC_130 NC_131 NC_132 NC_133 NC_134 NC_135 AT28HC256EPLCC32
.end
