.title KiCad schematic
U1 NC_01 NC_02 Net-_R3-Pad1_ Net-_R6-Pad1_ Net-_R4-Pad1_ Net-_R5-Pad1_ Net-_C5-Pad1_ GND VDDA Net-_R7-Pad2_ Net-_R8-Pad2_ Net-_R9-Pad2_ /GPIO1 /GPIO2 /GPIO3 NC_03 NC_04 NC_05 /OPTO1 /OPTO2 NC_06 NC_07 NC_08 VDD NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 VDD NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 Net-_1K1-Pad1_ NC_27 NC_28 NC_29 VDD STM32L433CCT6
SW1 GND Net-_C5-Pad1_ RST
C5 Net-_C5-Pad1_ GND 100nF
1K1 Net-_1K1-Pad1_ GND R1
T2 Net-_R11-Pad2_ NC_30 GND /OPTO1 TLP291
R10 VDD /OPTO1 1K
R11 NC_31 Net-_R11-Pad2_ 510
T1 Net-_R2-Pad2_ NC_32 GND /OPTO2 TLP291
R1 VDD /OPTO2 1K
R2 NC_33 Net-_R2-Pad2_ 510
T3 Net-_R12-Pad1_ GND NC_34 NC_35 TLP3556
R12 Net-_R12-Pad1_ NC_36 510
R7 NC_37 Net-_R7-Pad2_ 22
R8 NC_38 Net-_R8-Pad2_ 22
R9 NC_39 Net-_R9-Pad2_ 22
Y1 Net-_C1-Pad1_ NC_40 NC_41 Net-_C2-Pad1_ ABS25-32.768KHZ-6-T
C1 Net-_C1-Pad1_ GND 4.3pF
R3 Net-_R3-Pad1_ Net-_C1-Pad1_ 0R
C2 Net-_C2-Pad1_ GND 4.3pF
R6 Net-_R6-Pad1_ Net-_C2-Pad1_ 0R
X1 NC_42 NC_43 ABLS-8.000MHZ-B2-T
C4 Net-_C4-Pad1_ GND 20pF
R5 Net-_R5-Pad1_ Net-_C4-Pad1_ 0R
C3 Net-_C3-Pad1_ GND 20pF
R4 Net-_R4-Pad1_ Net-_C3-Pad1_ 0R
FB1 VDDA VDD 800mA 250m
C6 VDD GND 1uF
C7 VDD GND 100nF
C8 VDD GND 10nF
C9 VDDA GND 100nF
R13 /GPIO1 GND 10K
R14 /GPIO2 GND 10K
R15 /GPIO3 GND 10K
R16 NC_44 GND 10.1K
.end
