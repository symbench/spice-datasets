.title KiCad schematic
J1 -12V GND GND +12V Conn_01x04
J2 +12V +12V GND GND GND GND GND GND -12V -12V Conn_02x05_Odd_Even
J3 +12V +12V GND GND GND GND GND GND -12V -12V Conn_02x05_Odd_Even
J4 +12V +12V GND GND GND GND GND GND -12V -12V Conn_02x05_Odd_Even
J5 +12V +12V GND GND GND GND GND GND -12V -12V Conn_02x05_Odd_Even
J6 +12V +12V GND GND GND GND GND GND -12V -12V Conn_02x05_Odd_Even
C1 +12V GND 6800uF
C2 GND -12V 6800uF
R1 Net-_D1-Pad2_ +12V 1K
R2 -12V Net-_D2-Pad1_ 1K
D1 GND Net-_D1-Pad2_ +12V
D2 Net-_D2-Pad1_ GND -12V
H1 GND MountingHole_Pad
H2 GND MountingHole_Pad
H3 GND MountingHole_Pad
H4 GND MountingHole_Pad
J7 +12V +12V GND GND GND GND GND GND -12V -12V Conn_02x05_Odd_Even
.end
