.title KiCad schematic
U2 VCC GND /SCL /SDA NC_01 NC_02 NC_03 NC_04 GY-521
U1 VCC GND VCC Net-_C2-Pad1_ +3V3 MIC5219-3.3
C2 Net-_C2-Pad1_ GND 470p
C3 +3V3 GND 2.2uf
C1 VCC GND 2.2uf
R2 +3V3 /Temp 4.7k
R1 VCC Net-_R1-Pad2_ 47K
U4 GND /Temp VCC DS18B20
U3 NC_05 GND Net-_SW1-Pad3_ NC_06 NC_07 NC_08 TP4056-shield-6PIN
R3 Net-_R1-Pad2_ GND 10K
U6 Net-_C6-Pad1_ Net-_R1-Pad2_ /EN /RES /SCK /MISO /MOSI +3V3 GND /NSS /SCL /SDA /LED /Temp Net-_J2-Pad3_ Net-_J2-Pad2_ ESP-07S
D1 /RES Net-_C6-Pad1_ Schottky
R4 /EN +3V3 10K
R5 +3V3 Net-_C6-Pad1_ 10K
R6 GND /NSS 10K
C5 +3V3 GND 10uf
C4 +3V3 GND 100n
J1 /SDA GND PROG
U5 GND GND +3V3 /RES NC_09 NC_10 NC_11 NC_12 GND NC_13 NC_14 /SCK /MISO /MOSI /NSS GND LoRa_Ra-02
J2 GND Net-_J2-Pad2_ Net-_J2-Pad3_ /VCC_PROG PROG_con
SW1 /VCC_PROG VCC Net-_SW1-Pad3_ SW_SPDT
SW2 /VCC_PROG VCC Net-_SW1-Pad3_ SW_SPDT
SW3 Net-_C6-Pad1_ GND SW_Push
C6 Net-_C6-Pad1_ GND 100n
D2 /LED Net-_D2-Pad2_ LED
R7 +3V3 Net-_D2-Pad2_ 4.7k
C7 VCC GND 100n
.end
