.title KiCad schematic
R201 NC_01 NC_02 1k
R202 NC_03 NC_04 1k
R203 NC_05 NC_06 1k
R204 NC_07 NC_08 1k
R205 NC_09 NC_10 1k
R206 NC_11 NC_12 1k
R207 NC_13 NC_14 1k
R208 NC_15 NC_16 1k
.end
