.title KiCad schematic
R3 Net-_J3-Pad3_ Net-_J1-Pad1_ R
J1 Net-_J1-Pad1_ Net-_D1-Pad1_ 5V Sup
J3 Net-_J1-Pad1_ Net-_D1-Pad1_ Net-_J3-Pad3_ Net-_J3-Pad4_ Net-_J3-Pad5_ Net-_J3-Pad6_ Conn_01x06
J2 Net-_J2-Pad1_ Net-_J2-Pad2_ Net-_J1-Pad1_ Net-_D1-Pad1_ Conn_01x04
R2 Net-_R2-Pad1_ Net-_D2-Pad2_ R
D2 Net-_D1-Pad1_ Net-_D2-Pad2_ LED
D1 Net-_D1-Pad1_ Net-_D1-Pad2_ LED
R1 Net-_R1-Pad1_ Net-_D1-Pad2_ R
U1 Net-_J3-Pad3_ NC_01 NC_02 Net-_J2-Pad2_ Net-_J2-Pad1_ Net-_R1-Pad1_ Net-_J1-Pad1_ Net-_D1-Pad1_ Net-_R2-Pad1_ NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 Net-_J3-Pad4_ Net-_J3-Pad5_ Net-_J3-Pad6_ Net-_J1-Pad1_ NC_10 Net-_D1-Pad1_ NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 ATMEGA328P-PU
.end
