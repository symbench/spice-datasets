.title KiCad schematic
U8 /XBEE_VCC /TX_ISOLATED /RX_ISOLATED NC_01 NC_02 Net-_R21-Pad1_ NC_03 NC_04 GND NC_05 NC_06 NC_07 GND Net-_TP2-Pad1_ NC_08 NC_09 NC_10 NC_11 NC_12 XBP9B-DPST-001
C41 /XBEE_VCC GND 10uF
C40 /XBEE_VCC GND 0.01uF
U10 +3V3 GND CC_GPIO7 Net-_C44-Pad1_ Net-_R23-Pad2_ /XBEE_VCC TPS22918
R23 /XBEE_VCC Net-_R23-Pad2_ 0
C44 Net-_C44-Pad1_ GND 0.001uF
R24 CC_GPIO7 GND 100K
C46 GND +3V3 1uF
C42 /XBEE_VCC GND 22uF
TP2 Net-_TP2-Pad1_ Test_Point
R21 Net-_R21-Pad1_ Net-_D1-Pad2_ 330
D1 GND Net-_D1-Pad2_ LG L29K-F2J1-24-Z 
U9 /RX_ISOLATED GND +3V3 NC_13 NC_14 /XBEE_VCC /XBEE_VCC /TX_ISOLATED TXB0102DCU
C43 +3V3 GND 0.1uF
R22 /XBEE_VCC GND 100K
.end
