.title KiCad schematic
J1 +5V +5V -5V -5V +2V5 -2V5 GND GND +45V +45V GND GND -45V -45V GND GND /D_DATA /D_CLK /~D_CS /~D_RESET /~D_LOAD NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 PinDriverConnector
C5 +2V5 GND 100n
C6 -2V5 GND 100n
U1 +5V NC_20 NC_21 -2V5 +2V5 NC_22 NC_23 -5V GND /D_DATA /D_CLK /~D_CS NC_24 /~D_LOAD /~D_RESET +5V DAC7614U
C1 +5V GND 100n
C3 +5V GND 1u
C4 GND -5V 1u
C2 -5V GND 100n
.end
