.title KiCad schematic
X1 /RED /GREEN /BLUE NC_01 NC_02 GND GND GND NC_03 GND GND NC_04 Net-_R29-Pad2_ Net-_R30-Pad2_ NC_05 VGA
R42 NC_06 /RED 3.9K
R35 NC_07 /GREEN 3.9K
R31 NC_08 /BLUE 3.9K
R29 NC_09 Net-_R29-Pad2_ 82.5
R30 NC_10 Net-_R30-Pad2_ 82.5
R41 NC_11 /RED 2K
R36 NC_12 /GREEN 2K
R32 NC_13 /BLUE 2K
R40 NC_14 /RED 1K
R39 NC_15 /RED 510
R37 NC_16 /GREEN 1K
R38 NC_17 /GREEN 510
R33 NC_18 /BLUE 1K
R34 NC_19 /BLUE 510
.end
