.title KiCad schematic
J1 Net-_J1-Pad1_ Net-_J1-Pad2_ Net-_J1-Pad3_ NC_01 NC_02 GND RB1-125BAG1A
R1 Net-_R1-Pad1_ Net-_J1-Pad1_ 1k
R2 Net-_Q1-Pad2_ Net-_R1-Pad1_ 10k
U1 Net-_R1-Pad1_ Net-_J1-Pad2_ GND Net-_Q1-Pad2_ +9V LM7171
R4 +9V Net-_J1-Pad3_ 1k
Q1 Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_D1-Pad1_ 2N3904
R3 Net-_Q1-Pad1_ GND 450
D1 Net-_D1-Pad1_ +9V LTL2T3TBK5
BT1 +9V GND 9V
C1 +9V GND 33uF
C2 GND +9V C
Q2 Net-_J1-Pad3_ GND GND 2N3906
U2 GND Physical_Mount
U3 GND Physical_Mount
.end
