.title KiCad schematic
C15 +5V GND 0.1uF
J2 NC_01 NC_02 NC_03 NC_04 GND GND NC_05 NC_06 NC_07 NC_08 GND GND NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 IR_SIM_CLOCK NC_20 IR_SIM_RESET IR_SIM_IO RF_EN NC_21 MODE_SW NC_22 NC_23 NC_24 GND GND +5V +30V +5V +30V +5V 53885-0408
C6 SIM_VCC GND 1uF
U2 NC_25 NC_26 +5V NC_27 +5V NC_28 SIM_VCC SIM_IO SIM_RESET GND SIM_CLOCK NC_29 IR_SIM_CLOCK IR_SIM_RESET IR_SIM_IO NC_30 GND NCN4555MN
C5 +5V GND 0.1u
JP1 MODE_SW RF_EN SolderJumper_2_Open
R8 RF_EN GND 100k
C9 +8V GND 10uF
C2 Net-_C2-Pad1_ Net-_C2-Pad2_ 100pF
C1 Net-_C1-Pad1_ GND 33nF
R1 Net-_C3-Pad1_ Net-_C4-Pad1_ 12.1k
C3 Net-_C3-Pad1_ Net-_C3-Pad2_ 1.5nF
C4 Net-_C4-Pad1_ Net-_C3-Pad2_ 27nF
R3 Net-_C2-Pad1_ +8V 301k
C8 GND Net-_C8-Pad2_ 1uF
R4 Net-_C3-Pad1_ +30V 47.5k
R5 Net-_Q1-Pad4_ Net-_R5-Pad2_ 19.1
R6 Net-_Q1-Pad1_ Net-_C7-Pad1_ 1k
R7 Net-_Q1-Pad1_ GND 15m
C7 Net-_C7-Pad1_ GND 150pF
C10 +8V GND 470nF
R2 Net-_C3-Pad1_ GND 1.13k
C13 +30V GND 2.2uF
U1 Net-_C2-Pad2_ Net-_C1-Pad1_ NC_31 Net-_C3-Pad2_ Net-_C3-Pad1_ GND Net-_C7-Pad1_ Net-_R5-Pad2_ Net-_C8-Pad2_ +8V TPS40210DGQR
C16 +30V GND 0.1uF
C12 MODE_SW GND 1uF
C14 MODE_SW GND 10uF
C11 +30V GND +30V +30V GND GND 39uF
CR1 +30V Net-_CR1-Pad2_ B260-13-F
L1 Net-_CR1-Pad2_ +8V 24uH
J1 SIM_CLOCK SIM_RESET SIM_VCC SIM_IO NC_32 GND GND GND 47388-2001
Q1 Net-_Q1-Pad1_ Net-_Q1-Pad1_ Net-_Q1-Pad1_ Net-_Q1-Pad4_ Net-_CR1-Pad2_ Net-_CR1-Pad2_ Net-_CR1-Pad2_ Net-_CR1-Pad2_ Net-_CR1-Pad2_ CSD18543Q3AT
.end
