.title KiCad schematic
J1 /+12V_RAW /+12V_RAW GND GND GND GND GND GND /-12V_RAW /-12V_RAW EuroPower
R1 +12V /+12V_RAW 10R
R2 -12V /-12V_RAW 10R
C1 +12V GND 10uF
C2 GND -12V 10uF
U1 +12V GND +5V L7805
C3 +5V GND 10uF
J2 +5V +5V +12V +12V GND GND GND GND GND GND -12V -12V Interconnect
U2 +12V NC_01 +5V L7805
.end
