.title KiCad schematic
Q1 Net-_D1-Pad2_ Net-_F1-Pad1_ +24V Q_PMOS_GDS
R1 Net-_D1-Pad2_ GND R
D1 +24V Net-_D1-Pad2_ D_Zener
U1 +5V +5V +5V GND GND +24V +24V +5V +5V +5V GND GND +24V +24V +5V +5V +5V GND GND +24V +24V +5V +5V +5V GND GND GND GND GND GND GND Net-_U1-Pad5F_ Net-_U1-Pad5F_ GND GND GND GND GND GND GND NC_01 GND GND GND GND GND NC_02 Net-_R3-Pad2_ Net-_R2-Pad2_ LTM8022or8023
R2 GND Net-_R2-Pad2_ R
R3 GND Net-_R3-Pad2_ R
C4 +5V GND C
C3 +5V GND CP
C2 +24V GND CP
C1 +24V GND C
U2 +3V3 +3V3 +3V3 GND GND +24V +24V +3V3 +3V3 +3V3 GND GND +24V +24V +3V3 +3V3 +3V3 GND GND +24V +24V +3V3 +3V3 +3V3 GND GND GND GND GND GND GND Net-_U2-Pad5F_ Net-_U2-Pad5F_ GND GND GND GND GND GND GND NC_03 GND GND GND GND GND NC_04 Net-_R5-Pad2_ Net-_R4-Pad2_ LTM8022or8023
R4 GND Net-_R4-Pad2_ R
R5 GND Net-_R5-Pad2_ R
C8 +3V3 GND C
C7 +3V3 GND CP
C6 +24V GND CP
C5 +24V GND C
F1 Net-_F1-Pad1_ +BATT Fuse
D2 +24V GND D_Zener
D3 +24V GND D_Zener
D4 +5V GND D_Zener
D5 +5V GND D_Zener
D6 +3V3 GND D_Zener
D7 +3V3 GND D_Zener
.end
