.title KiCad schematic
U1 NC_01 Net-_U1-Pad2_ Net-_U1-Pad2_ NC_02 MINI-360
U3 Net-_U3-Pad1_ NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 Net-_U3-Pad1_ NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 Net-_U3-Pad38_ Net-_U3-Pad38_ ESP32-WROOM
.end
